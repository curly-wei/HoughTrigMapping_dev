library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
 
entity UT3_0_SL6 is
 
Port (
           SL6_row1  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row2  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row3  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row4  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row5  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row6  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row7  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row8  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row9  : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row10 : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row11 : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row12 : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row13 : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row14 : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row15 : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_row16 : out  STD_LOGIC_VECTOR (79 downto 40);
           SL6_TS    : in   STD_LOGIC_VECTOR (160 downto 0));
end UT3_0_SL6;
 
 
architecture Behavioral of UT3_0_SL6 is
 
begin
 
SL6_row1(40)<=SL6_TS(28) or SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) ;
SL6_row1(41)<=SL6_TS(30) or SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) ;
SL6_row1(42)<=SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) ;
SL6_row1(43)<=SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) ;
SL6_row1(44)<=SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) ;
SL6_row1(45)<=SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) ;
SL6_row1(46)<=SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) ;
SL6_row1(47)<=SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) ;
SL6_row1(48)<=SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) ;
SL6_row1(49)<=SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) ;
SL6_row1(50)<=SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) ;
SL6_row1(51)<=SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) ;
SL6_row1(52)<=SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) ;
SL6_row1(53)<=SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) ;
SL6_row1(54)<=SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) ;
SL6_row1(55)<=SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) ;
SL6_row1(56)<=SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) ;
SL6_row1(57)<=SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) ;
SL6_row1(58)<=SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) ;
SL6_row1(59)<=SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) ;
SL6_row1(60)<=SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) ;
SL6_row1(61)<=SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) ;
SL6_row1(62)<=SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) ;
SL6_row1(63)<=SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) ;
SL6_row1(64)<=SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) ;
SL6_row1(65)<=SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) ;
SL6_row1(66)<=SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) ;
SL6_row1(67)<=SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) ;
SL6_row1(68)<=SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) ;
SL6_row1(69)<=SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) ;
SL6_row1(70)<=SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) ;
SL6_row1(71)<=SL6_TS(90) or SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) or SL6_TS(97) or SL6_TS(98) ;
SL6_row1(72)<=SL6_TS(92) or SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) or SL6_TS(97) or SL6_TS(98) or SL6_TS(99) or SL6_TS(100) ;
SL6_row1(73)<=SL6_TS(94) or SL6_TS(95) or SL6_TS(96) or SL6_TS(97) or SL6_TS(98) or SL6_TS(99) or SL6_TS(100) or SL6_TS(101) or SL6_TS(102) ;
SL6_row1(74)<=SL6_TS(96) or SL6_TS(97) or SL6_TS(98) or SL6_TS(99) or SL6_TS(100) or SL6_TS(101) or SL6_TS(102) or SL6_TS(103) or SL6_TS(104) ;
SL6_row1(75)<=SL6_TS(98) or SL6_TS(99) or SL6_TS(100) or SL6_TS(101) or SL6_TS(102) or SL6_TS(103) or SL6_TS(104) or SL6_TS(105) or SL6_TS(106) ;
SL6_row1(76)<=SL6_TS(100) or SL6_TS(101) or SL6_TS(102) or SL6_TS(103) or SL6_TS(104) or SL6_TS(105) or SL6_TS(106) or SL6_TS(107) or SL6_TS(108) ;
SL6_row1(77)<=SL6_TS(102) or SL6_TS(103) or SL6_TS(104) or SL6_TS(105) or SL6_TS(106) or SL6_TS(107) or SL6_TS(108) or SL6_TS(109) or SL6_TS(110) ;
SL6_row1(78)<=SL6_TS(104) or SL6_TS(105) or SL6_TS(106) or SL6_TS(107) or SL6_TS(108) or SL6_TS(109) or SL6_TS(110) or SL6_TS(111) or SL6_TS(112) ;
SL6_row1(79)<=SL6_TS(106) or SL6_TS(107) or SL6_TS(108) or SL6_TS(109) or SL6_TS(110) or SL6_TS(111) or SL6_TS(112) or SL6_TS(113) or SL6_TS(114) ;
SL6_row2(40)<=SL6_TS(23) or SL6_TS(24) or SL6_TS(25) or SL6_TS(26) or SL6_TS(27) or SL6_TS(28) or SL6_TS(29) ;
SL6_row2(41)<=SL6_TS(25) or SL6_TS(26) or SL6_TS(27) or SL6_TS(28) or SL6_TS(29) or SL6_TS(30) or SL6_TS(31) ;
SL6_row2(42)<=SL6_TS(27) or SL6_TS(28) or SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) or SL6_TS(33) ;
SL6_row2(43)<=SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) ;
SL6_row2(44)<=SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) ;
SL6_row2(45)<=SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) ;
SL6_row2(46)<=SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) ;
SL6_row2(47)<=SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) ;
SL6_row2(48)<=SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) ;
SL6_row2(49)<=SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) ;
SL6_row2(50)<=SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) ;
SL6_row2(51)<=SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) ;
SL6_row2(52)<=SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) ;
SL6_row2(53)<=SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) ;
SL6_row2(54)<=SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) ;
SL6_row2(55)<=SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) ;
SL6_row2(56)<=SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) ;
SL6_row2(57)<=SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) ;
SL6_row2(58)<=SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) ;
SL6_row2(59)<=SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) ;
SL6_row2(60)<=SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) ;
SL6_row2(61)<=SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) ;
SL6_row2(62)<=SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) ;
SL6_row2(63)<=SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) ;
SL6_row2(64)<=SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) ;
SL6_row2(65)<=SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) ;
SL6_row2(66)<=SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) ;
SL6_row2(67)<=SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) ;
SL6_row2(68)<=SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) ;
SL6_row2(69)<=SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) ;
SL6_row2(70)<=SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) ;
SL6_row2(71)<=SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) ;
SL6_row2(72)<=SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) or SL6_TS(93) ;
SL6_row2(73)<=SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) or SL6_TS(95) ;
SL6_row2(74)<=SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) or SL6_TS(97) ;
SL6_row2(75)<=SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) or SL6_TS(97) or SL6_TS(98) or SL6_TS(99) ;
SL6_row2(76)<=SL6_TS(95) or SL6_TS(96) or SL6_TS(97) or SL6_TS(98) or SL6_TS(99) or SL6_TS(100) or SL6_TS(101) ;
SL6_row2(77)<=SL6_TS(97) or SL6_TS(98) or SL6_TS(99) or SL6_TS(100) or SL6_TS(101) or SL6_TS(102) or SL6_TS(103) ;
SL6_row2(78)<=SL6_TS(99) or SL6_TS(100) or SL6_TS(101) or SL6_TS(102) or SL6_TS(103) or SL6_TS(104) or SL6_TS(105) ;
SL6_row2(79)<=SL6_TS(101) or SL6_TS(102) or SL6_TS(103) or SL6_TS(104) or SL6_TS(105) or SL6_TS(106) or SL6_TS(107) ;
SL6_row3(40)<=SL6_TS(19) or SL6_TS(20) or SL6_TS(21) or SL6_TS(22) or SL6_TS(23) or SL6_TS(24) ;
SL6_row3(41)<=SL6_TS(21) or SL6_TS(22) or SL6_TS(23) or SL6_TS(24) or SL6_TS(25) or SL6_TS(26) ;
SL6_row3(42)<=SL6_TS(23) or SL6_TS(24) or SL6_TS(25) or SL6_TS(26) or SL6_TS(27) or SL6_TS(28) ;
SL6_row3(43)<=SL6_TS(25) or SL6_TS(26) or SL6_TS(27) or SL6_TS(28) or SL6_TS(29) or SL6_TS(30) ;
SL6_row3(44)<=SL6_TS(27) or SL6_TS(28) or SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) ;
SL6_row3(45)<=SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) ;
SL6_row3(46)<=SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) ;
SL6_row3(47)<=SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) ;
SL6_row3(48)<=SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) ;
SL6_row3(49)<=SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) ;
SL6_row3(50)<=SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) ;
SL6_row3(51)<=SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) ;
SL6_row3(52)<=SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) ;
SL6_row3(53)<=SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) ;
SL6_row3(54)<=SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) ;
SL6_row3(55)<=SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) ;
SL6_row3(56)<=SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) ;
SL6_row3(57)<=SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) ;
SL6_row3(58)<=SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) ;
SL6_row3(59)<=SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) ;
SL6_row3(60)<=SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) ;
SL6_row3(61)<=SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) ;
SL6_row3(62)<=SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) ;
SL6_row3(63)<=SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) ;
SL6_row3(64)<=SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) ;
SL6_row3(65)<=SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) ;
SL6_row3(66)<=SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) ;
SL6_row3(67)<=SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) ;
SL6_row3(68)<=SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) ;
SL6_row3(69)<=SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) ;
SL6_row3(70)<=SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) ;
SL6_row3(71)<=SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) ;
SL6_row3(72)<=SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) ;
SL6_row3(73)<=SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) ;
SL6_row3(74)<=SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) ;
SL6_row3(75)<=SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) ;
SL6_row3(76)<=SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) ;
SL6_row3(77)<=SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) or SL6_TS(97) or SL6_TS(98) ;
SL6_row3(78)<=SL6_TS(95) or SL6_TS(96) or SL6_TS(97) or SL6_TS(98) or SL6_TS(99) or SL6_TS(100) ;
SL6_row3(79)<=SL6_TS(97) or SL6_TS(98) or SL6_TS(99) or SL6_TS(100) or SL6_TS(101) or SL6_TS(102) ;
SL6_row4(40)<=SL6_TS(15) or SL6_TS(16) or SL6_TS(17) or SL6_TS(18) or SL6_TS(19) or SL6_TS(20) ;
SL6_row4(41)<=SL6_TS(17) or SL6_TS(18) or SL6_TS(19) or SL6_TS(20) or SL6_TS(21) or SL6_TS(22) ;
SL6_row4(42)<=SL6_TS(19) or SL6_TS(20) or SL6_TS(21) or SL6_TS(22) or SL6_TS(23) or SL6_TS(24) ;
SL6_row4(43)<=SL6_TS(21) or SL6_TS(22) or SL6_TS(23) or SL6_TS(24) or SL6_TS(25) or SL6_TS(26) ;
SL6_row4(44)<=SL6_TS(23) or SL6_TS(24) or SL6_TS(25) or SL6_TS(26) or SL6_TS(27) or SL6_TS(28) ;
SL6_row4(45)<=SL6_TS(25) or SL6_TS(26) or SL6_TS(27) or SL6_TS(28) or SL6_TS(29) or SL6_TS(30) ;
SL6_row4(46)<=SL6_TS(27) or SL6_TS(28) or SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) ;
SL6_row4(47)<=SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) ;
SL6_row4(48)<=SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) ;
SL6_row4(49)<=SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) ;
SL6_row4(50)<=SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) ;
SL6_row4(51)<=SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) ;
SL6_row4(52)<=SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) ;
SL6_row4(53)<=SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) ;
SL6_row4(54)<=SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) ;
SL6_row4(55)<=SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) ;
SL6_row4(56)<=SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) ;
SL6_row4(57)<=SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) ;
SL6_row4(58)<=SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) ;
SL6_row4(59)<=SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) ;
SL6_row4(60)<=SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) ;
SL6_row4(61)<=SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) ;
SL6_row4(62)<=SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) ;
SL6_row4(63)<=SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) ;
SL6_row4(64)<=SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) ;
SL6_row4(65)<=SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) ;
SL6_row4(66)<=SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) ;
SL6_row4(67)<=SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) ;
SL6_row4(68)<=SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) ;
SL6_row4(69)<=SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) ;
SL6_row4(70)<=SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) ;
SL6_row4(71)<=SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) ;
SL6_row4(72)<=SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) ;
SL6_row4(73)<=SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) ;
SL6_row4(74)<=SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) ;
SL6_row4(75)<=SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) ;
SL6_row4(76)<=SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) ;
SL6_row4(77)<=SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) ;
SL6_row4(78)<=SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) ;
SL6_row4(79)<=SL6_TS(93) or SL6_TS(94) or SL6_TS(95) or SL6_TS(96) or SL6_TS(97) or SL6_TS(98) ;
SL6_row5(40)<=SL6_TS(12) or SL6_TS(13) or SL6_TS(14) or SL6_TS(15) or SL6_TS(16) ;
SL6_row5(41)<=SL6_TS(14) or SL6_TS(15) or SL6_TS(16) or SL6_TS(17) or SL6_TS(18) ;
SL6_row5(42)<=SL6_TS(16) or SL6_TS(17) or SL6_TS(18) or SL6_TS(19) or SL6_TS(20) ;
SL6_row5(43)<=SL6_TS(18) or SL6_TS(19) or SL6_TS(20) or SL6_TS(21) or SL6_TS(22) ;
SL6_row5(44)<=SL6_TS(20) or SL6_TS(21) or SL6_TS(22) or SL6_TS(23) or SL6_TS(24) ;
SL6_row5(45)<=SL6_TS(22) or SL6_TS(23) or SL6_TS(24) or SL6_TS(25) or SL6_TS(26) ;
SL6_row5(46)<=SL6_TS(24) or SL6_TS(25) or SL6_TS(26) or SL6_TS(27) or SL6_TS(28) ;
SL6_row5(47)<=SL6_TS(26) or SL6_TS(27) or SL6_TS(28) or SL6_TS(29) or SL6_TS(30) ;
SL6_row5(48)<=SL6_TS(28) or SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) ;
SL6_row5(49)<=SL6_TS(30) or SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) ;
SL6_row5(50)<=SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) ;
SL6_row5(51)<=SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) ;
SL6_row5(52)<=SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) ;
SL6_row5(53)<=SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) ;
SL6_row5(54)<=SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) ;
SL6_row5(55)<=SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) ;
SL6_row5(56)<=SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) ;
SL6_row5(57)<=SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) ;
SL6_row5(58)<=SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) ;
SL6_row5(59)<=SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) ;
SL6_row5(60)<=SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) ;
SL6_row5(61)<=SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) ;
SL6_row5(62)<=SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) ;
SL6_row5(63)<=SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) ;
SL6_row5(64)<=SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) ;
SL6_row5(65)<=SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) ;
SL6_row5(66)<=SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) ;
SL6_row5(67)<=SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) ;
SL6_row5(68)<=SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) ;
SL6_row5(69)<=SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) ;
SL6_row5(70)<=SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) ;
SL6_row5(71)<=SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) ;
SL6_row5(72)<=SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) ;
SL6_row5(73)<=SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) ;
SL6_row5(74)<=SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) ;
SL6_row5(75)<=SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) ;
SL6_row5(76)<=SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) ;
SL6_row5(77)<=SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) or SL6_TS(90) ;
SL6_row5(78)<=SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) or SL6_TS(92) ;
SL6_row5(79)<=SL6_TS(90) or SL6_TS(91) or SL6_TS(92) or SL6_TS(93) or SL6_TS(94) ;
SL6_row6(40)<=SL6_TS(10) or SL6_TS(11) or SL6_TS(12) or SL6_TS(13) ;
SL6_row6(41)<=SL6_TS(12) or SL6_TS(13) or SL6_TS(14) or SL6_TS(15) ;
SL6_row6(42)<=SL6_TS(14) or SL6_TS(15) or SL6_TS(16) or SL6_TS(17) ;
SL6_row6(43)<=SL6_TS(16) or SL6_TS(17) or SL6_TS(18) or SL6_TS(19) ;
SL6_row6(44)<=SL6_TS(18) or SL6_TS(19) or SL6_TS(20) or SL6_TS(21) ;
SL6_row6(45)<=SL6_TS(20) or SL6_TS(21) or SL6_TS(22) or SL6_TS(23) ;
SL6_row6(46)<=SL6_TS(22) or SL6_TS(23) or SL6_TS(24) or SL6_TS(25) ;
SL6_row6(47)<=SL6_TS(24) or SL6_TS(25) or SL6_TS(26) or SL6_TS(27) ;
SL6_row6(48)<=SL6_TS(26) or SL6_TS(27) or SL6_TS(28) or SL6_TS(29) ;
SL6_row6(49)<=SL6_TS(28) or SL6_TS(29) or SL6_TS(30) or SL6_TS(31) ;
SL6_row6(50)<=SL6_TS(30) or SL6_TS(31) or SL6_TS(32) or SL6_TS(33) ;
SL6_row6(51)<=SL6_TS(32) or SL6_TS(33) or SL6_TS(34) or SL6_TS(35) ;
SL6_row6(52)<=SL6_TS(34) or SL6_TS(35) or SL6_TS(36) or SL6_TS(37) ;
SL6_row6(53)<=SL6_TS(36) or SL6_TS(37) or SL6_TS(38) or SL6_TS(39) ;
SL6_row6(54)<=SL6_TS(38) or SL6_TS(39) or SL6_TS(40) or SL6_TS(41) ;
SL6_row6(55)<=SL6_TS(40) or SL6_TS(41) or SL6_TS(42) or SL6_TS(43) ;
SL6_row6(56)<=SL6_TS(42) or SL6_TS(43) or SL6_TS(44) or SL6_TS(45) ;
SL6_row6(57)<=SL6_TS(44) or SL6_TS(45) or SL6_TS(46) or SL6_TS(47) ;
SL6_row6(58)<=SL6_TS(46) or SL6_TS(47) or SL6_TS(48) or SL6_TS(49) ;
SL6_row6(59)<=SL6_TS(48) or SL6_TS(49) or SL6_TS(50) or SL6_TS(51) ;
SL6_row6(60)<=SL6_TS(50) or SL6_TS(51) or SL6_TS(52) or SL6_TS(53) ;
SL6_row6(61)<=SL6_TS(52) or SL6_TS(53) or SL6_TS(54) or SL6_TS(55) ;
SL6_row6(62)<=SL6_TS(54) or SL6_TS(55) or SL6_TS(56) or SL6_TS(57) ;
SL6_row6(63)<=SL6_TS(56) or SL6_TS(57) or SL6_TS(58) or SL6_TS(59) ;
SL6_row6(64)<=SL6_TS(58) or SL6_TS(59) or SL6_TS(60) or SL6_TS(61) ;
SL6_row6(65)<=SL6_TS(60) or SL6_TS(61) or SL6_TS(62) or SL6_TS(63) ;
SL6_row6(66)<=SL6_TS(62) or SL6_TS(63) or SL6_TS(64) or SL6_TS(65) ;
SL6_row6(67)<=SL6_TS(64) or SL6_TS(65) or SL6_TS(66) or SL6_TS(67) ;
SL6_row6(68)<=SL6_TS(66) or SL6_TS(67) or SL6_TS(68) or SL6_TS(69) ;
SL6_row6(69)<=SL6_TS(68) or SL6_TS(69) or SL6_TS(70) or SL6_TS(71) ;
SL6_row6(70)<=SL6_TS(70) or SL6_TS(71) or SL6_TS(72) or SL6_TS(73) ;
SL6_row6(71)<=SL6_TS(72) or SL6_TS(73) or SL6_TS(74) or SL6_TS(75) ;
SL6_row6(72)<=SL6_TS(74) or SL6_TS(75) or SL6_TS(76) or SL6_TS(77) ;
SL6_row6(73)<=SL6_TS(76) or SL6_TS(77) or SL6_TS(78) or SL6_TS(79) ;
SL6_row6(74)<=SL6_TS(78) or SL6_TS(79) or SL6_TS(80) or SL6_TS(81) ;
SL6_row6(75)<=SL6_TS(80) or SL6_TS(81) or SL6_TS(82) or SL6_TS(83) ;
SL6_row6(76)<=SL6_TS(82) or SL6_TS(83) or SL6_TS(84) or SL6_TS(85) ;
SL6_row6(77)<=SL6_TS(84) or SL6_TS(85) or SL6_TS(86) or SL6_TS(87) ;
SL6_row6(78)<=SL6_TS(86) or SL6_TS(87) or SL6_TS(88) or SL6_TS(89) ;
SL6_row6(79)<=SL6_TS(88) or SL6_TS(89) or SL6_TS(90) or SL6_TS(91) ;
SL6_row7(40)<=SL6_TS(9) or SL6_TS(10) or SL6_TS(11) ;
SL6_row7(41)<=SL6_TS(11) or SL6_TS(12) or SL6_TS(13) ;
SL6_row7(42)<=SL6_TS(13) or SL6_TS(14) or SL6_TS(15) ;
SL6_row7(43)<=SL6_TS(15) or SL6_TS(16) or SL6_TS(17) ;
SL6_row7(44)<=SL6_TS(17) or SL6_TS(18) or SL6_TS(19) ;
SL6_row7(45)<=SL6_TS(19) or SL6_TS(20) or SL6_TS(21) ;
SL6_row7(46)<=SL6_TS(21) or SL6_TS(22) or SL6_TS(23) ;
SL6_row7(47)<=SL6_TS(23) or SL6_TS(24) or SL6_TS(25) ;
SL6_row7(48)<=SL6_TS(25) or SL6_TS(26) or SL6_TS(27) ;
SL6_row7(49)<=SL6_TS(27) or SL6_TS(28) or SL6_TS(29) ;
SL6_row7(50)<=SL6_TS(29) or SL6_TS(30) or SL6_TS(31) ;
SL6_row7(51)<=SL6_TS(31) or SL6_TS(32) or SL6_TS(33) ;
SL6_row7(52)<=SL6_TS(33) or SL6_TS(34) or SL6_TS(35) ;
SL6_row7(53)<=SL6_TS(35) or SL6_TS(36) or SL6_TS(37) ;
SL6_row7(54)<=SL6_TS(37) or SL6_TS(38) or SL6_TS(39) ;
SL6_row7(55)<=SL6_TS(39) or SL6_TS(40) or SL6_TS(41) ;
SL6_row7(56)<=SL6_TS(41) or SL6_TS(42) or SL6_TS(43) ;
SL6_row7(57)<=SL6_TS(43) or SL6_TS(44) or SL6_TS(45) ;
SL6_row7(58)<=SL6_TS(45) or SL6_TS(46) or SL6_TS(47) ;
SL6_row7(59)<=SL6_TS(47) or SL6_TS(48) or SL6_TS(49) ;
SL6_row7(60)<=SL6_TS(49) or SL6_TS(50) or SL6_TS(51) ;
SL6_row7(61)<=SL6_TS(51) or SL6_TS(52) or SL6_TS(53) ;
SL6_row7(62)<=SL6_TS(53) or SL6_TS(54) or SL6_TS(55) ;
SL6_row7(63)<=SL6_TS(55) or SL6_TS(56) or SL6_TS(57) ;
SL6_row7(64)<=SL6_TS(57) or SL6_TS(58) or SL6_TS(59) ;
SL6_row7(65)<=SL6_TS(59) or SL6_TS(60) or SL6_TS(61) ;
SL6_row7(66)<=SL6_TS(61) or SL6_TS(62) or SL6_TS(63) ;
SL6_row7(67)<=SL6_TS(63) or SL6_TS(64) or SL6_TS(65) ;
SL6_row7(68)<=SL6_TS(65) or SL6_TS(66) or SL6_TS(67) ;
SL6_row7(69)<=SL6_TS(67) or SL6_TS(68) or SL6_TS(69) ;
SL6_row7(70)<=SL6_TS(69) or SL6_TS(70) or SL6_TS(71) ;
SL6_row7(71)<=SL6_TS(71) or SL6_TS(72) or SL6_TS(73) ;
SL6_row7(72)<=SL6_TS(73) or SL6_TS(74) or SL6_TS(75) ;
SL6_row7(73)<=SL6_TS(75) or SL6_TS(76) or SL6_TS(77) ;
SL6_row7(74)<=SL6_TS(77) or SL6_TS(78) or SL6_TS(79) ;
SL6_row7(75)<=SL6_TS(79) or SL6_TS(80) or SL6_TS(81) ;
SL6_row7(76)<=SL6_TS(81) or SL6_TS(82) or SL6_TS(83) ;
SL6_row7(77)<=SL6_TS(83) or SL6_TS(84) or SL6_TS(85) ;
SL6_row7(78)<=SL6_TS(85) or SL6_TS(86) or SL6_TS(87) ;
SL6_row7(79)<=SL6_TS(87) or SL6_TS(88) or SL6_TS(89) ;
SL6_row8(40)<=SL6_TS(7) or SL6_TS(8) or SL6_TS(9) or SL6_TS(10) ;
SL6_row8(41)<=SL6_TS(9) or SL6_TS(10) or SL6_TS(11) or SL6_TS(12) ;
SL6_row8(42)<=SL6_TS(11) or SL6_TS(12) or SL6_TS(13) or SL6_TS(14) ;
SL6_row8(43)<=SL6_TS(13) or SL6_TS(14) or SL6_TS(15) or SL6_TS(16) ;
SL6_row8(44)<=SL6_TS(15) or SL6_TS(16) or SL6_TS(17) or SL6_TS(18) ;
SL6_row8(45)<=SL6_TS(17) or SL6_TS(18) or SL6_TS(19) or SL6_TS(20) ;
SL6_row8(46)<=SL6_TS(19) or SL6_TS(20) or SL6_TS(21) or SL6_TS(22) ;
SL6_row8(47)<=SL6_TS(21) or SL6_TS(22) or SL6_TS(23) or SL6_TS(24) ;
SL6_row8(48)<=SL6_TS(23) or SL6_TS(24) or SL6_TS(25) or SL6_TS(26) ;
SL6_row8(49)<=SL6_TS(25) or SL6_TS(26) or SL6_TS(27) or SL6_TS(28) ;
SL6_row8(50)<=SL6_TS(27) or SL6_TS(28) or SL6_TS(29) or SL6_TS(30) ;
SL6_row8(51)<=SL6_TS(29) or SL6_TS(30) or SL6_TS(31) or SL6_TS(32) ;
SL6_row8(52)<=SL6_TS(31) or SL6_TS(32) or SL6_TS(33) or SL6_TS(34) ;
SL6_row8(53)<=SL6_TS(33) or SL6_TS(34) or SL6_TS(35) or SL6_TS(36) ;
SL6_row8(54)<=SL6_TS(35) or SL6_TS(36) or SL6_TS(37) or SL6_TS(38) ;
SL6_row8(55)<=SL6_TS(37) or SL6_TS(38) or SL6_TS(39) or SL6_TS(40) ;
SL6_row8(56)<=SL6_TS(39) or SL6_TS(40) or SL6_TS(41) or SL6_TS(42) ;
SL6_row8(57)<=SL6_TS(41) or SL6_TS(42) or SL6_TS(43) or SL6_TS(44) ;
SL6_row8(58)<=SL6_TS(43) or SL6_TS(44) or SL6_TS(45) or SL6_TS(46) ;
SL6_row8(59)<=SL6_TS(45) or SL6_TS(46) or SL6_TS(47) or SL6_TS(48) ;
SL6_row8(60)<=SL6_TS(47) or SL6_TS(48) or SL6_TS(49) or SL6_TS(50) ;
SL6_row8(61)<=SL6_TS(49) or SL6_TS(50) or SL6_TS(51) or SL6_TS(52) ;
SL6_row8(62)<=SL6_TS(51) or SL6_TS(52) or SL6_TS(53) or SL6_TS(54) ;
SL6_row8(63)<=SL6_TS(53) or SL6_TS(54) or SL6_TS(55) or SL6_TS(56) ;
SL6_row8(64)<=SL6_TS(55) or SL6_TS(56) or SL6_TS(57) or SL6_TS(58) ;
SL6_row8(65)<=SL6_TS(57) or SL6_TS(58) or SL6_TS(59) or SL6_TS(60) ;
SL6_row8(66)<=SL6_TS(59) or SL6_TS(60) or SL6_TS(61) or SL6_TS(62) ;
SL6_row8(67)<=SL6_TS(61) or SL6_TS(62) or SL6_TS(63) or SL6_TS(64) ;
SL6_row8(68)<=SL6_TS(63) or SL6_TS(64) or SL6_TS(65) or SL6_TS(66) ;
SL6_row8(69)<=SL6_TS(65) or SL6_TS(66) or SL6_TS(67) or SL6_TS(68) ;
SL6_row8(70)<=SL6_TS(67) or SL6_TS(68) or SL6_TS(69) or SL6_TS(70) ;
SL6_row8(71)<=SL6_TS(69) or SL6_TS(70) or SL6_TS(71) or SL6_TS(72) ;
SL6_row8(72)<=SL6_TS(71) or SL6_TS(72) or SL6_TS(73) or SL6_TS(74) ;
SL6_row8(73)<=SL6_TS(73) or SL6_TS(74) or SL6_TS(75) or SL6_TS(76) ;
SL6_row8(74)<=SL6_TS(75) or SL6_TS(76) or SL6_TS(77) or SL6_TS(78) ;
SL6_row8(75)<=SL6_TS(77) or SL6_TS(78) or SL6_TS(79) or SL6_TS(80) ;
SL6_row8(76)<=SL6_TS(79) or SL6_TS(80) or SL6_TS(81) or SL6_TS(82) ;
SL6_row8(77)<=SL6_TS(81) or SL6_TS(82) or SL6_TS(83) or SL6_TS(84) ;
SL6_row8(78)<=SL6_TS(83) or SL6_TS(84) or SL6_TS(85) or SL6_TS(86) ;
SL6_row8(79)<=SL6_TS(85) or SL6_TS(86) or SL6_TS(87) or SL6_TS(88) ;
SL6_row9(40)<=SL6_TS(6) or SL6_TS(7) or SL6_TS(8) ;
SL6_row9(41)<=SL6_TS(8) or SL6_TS(9) or SL6_TS(10) ;
SL6_row9(42)<=SL6_TS(10) or SL6_TS(11) or SL6_TS(12) ;
SL6_row9(43)<=SL6_TS(12) or SL6_TS(13) or SL6_TS(14) ;
SL6_row9(44)<=SL6_TS(14) or SL6_TS(15) or SL6_TS(16) ;
SL6_row9(45)<=SL6_TS(16) or SL6_TS(17) or SL6_TS(18) ;
SL6_row9(46)<=SL6_TS(18) or SL6_TS(19) or SL6_TS(20) ;
SL6_row9(47)<=SL6_TS(20) or SL6_TS(21) or SL6_TS(22) ;
SL6_row9(48)<=SL6_TS(22) or SL6_TS(23) or SL6_TS(24) ;
SL6_row9(49)<=SL6_TS(24) or SL6_TS(25) or SL6_TS(26) ;
SL6_row9(50)<=SL6_TS(26) or SL6_TS(27) or SL6_TS(28) ;
SL6_row9(51)<=SL6_TS(28) or SL6_TS(29) or SL6_TS(30) ;
SL6_row9(52)<=SL6_TS(30) or SL6_TS(31) or SL6_TS(32) ;
SL6_row9(53)<=SL6_TS(32) or SL6_TS(33) or SL6_TS(34) ;
SL6_row9(54)<=SL6_TS(34) or SL6_TS(35) or SL6_TS(36) ;
SL6_row9(55)<=SL6_TS(36) or SL6_TS(37) or SL6_TS(38) ;
SL6_row9(56)<=SL6_TS(38) or SL6_TS(39) or SL6_TS(40) ;
SL6_row9(57)<=SL6_TS(40) or SL6_TS(41) or SL6_TS(42) ;
SL6_row9(58)<=SL6_TS(42) or SL6_TS(43) or SL6_TS(44) ;
SL6_row9(59)<=SL6_TS(44) or SL6_TS(45) or SL6_TS(46) ;
SL6_row9(60)<=SL6_TS(46) or SL6_TS(47) or SL6_TS(48) ;
SL6_row9(61)<=SL6_TS(48) or SL6_TS(49) or SL6_TS(50) ;
SL6_row9(62)<=SL6_TS(50) or SL6_TS(51) or SL6_TS(52) ;
SL6_row9(63)<=SL6_TS(52) or SL6_TS(53) or SL6_TS(54) ;
SL6_row9(64)<=SL6_TS(54) or SL6_TS(55) or SL6_TS(56) ;
SL6_row9(65)<=SL6_TS(56) or SL6_TS(57) or SL6_TS(58) ;
SL6_row9(66)<=SL6_TS(58) or SL6_TS(59) or SL6_TS(60) ;
SL6_row9(67)<=SL6_TS(60) or SL6_TS(61) or SL6_TS(62) ;
SL6_row9(68)<=SL6_TS(62) or SL6_TS(63) or SL6_TS(64) ;
SL6_row9(69)<=SL6_TS(64) or SL6_TS(65) or SL6_TS(66) ;
SL6_row9(70)<=SL6_TS(66) or SL6_TS(67) or SL6_TS(68) ;
SL6_row9(71)<=SL6_TS(68) or SL6_TS(69) or SL6_TS(70) ;
SL6_row9(72)<=SL6_TS(70) or SL6_TS(71) or SL6_TS(72) ;
SL6_row9(73)<=SL6_TS(72) or SL6_TS(73) or SL6_TS(74) ;
SL6_row9(74)<=SL6_TS(74) or SL6_TS(75) or SL6_TS(76) ;
SL6_row9(75)<=SL6_TS(76) or SL6_TS(77) or SL6_TS(78) ;
SL6_row9(76)<=SL6_TS(78) or SL6_TS(79) or SL6_TS(80) ;
SL6_row9(77)<=SL6_TS(80) or SL6_TS(81) or SL6_TS(82) ;
SL6_row9(78)<=SL6_TS(82) or SL6_TS(83) or SL6_TS(84) ;
SL6_row9(79)<=SL6_TS(84) or SL6_TS(85) or SL6_TS(86) ;
SL6_row10(40)<=SL6_TS(5) or SL6_TS(6) or SL6_TS(7) ;
SL6_row10(41)<=SL6_TS(7) or SL6_TS(8) or SL6_TS(9) ;
SL6_row10(42)<=SL6_TS(9) or SL6_TS(10) or SL6_TS(11) ;
SL6_row10(43)<=SL6_TS(11) or SL6_TS(12) or SL6_TS(13) ;
SL6_row10(44)<=SL6_TS(13) or SL6_TS(14) or SL6_TS(15) ;
SL6_row10(45)<=SL6_TS(15) or SL6_TS(16) or SL6_TS(17) ;
SL6_row10(46)<=SL6_TS(17) or SL6_TS(18) or SL6_TS(19) ;
SL6_row10(47)<=SL6_TS(19) or SL6_TS(20) or SL6_TS(21) ;
SL6_row10(48)<=SL6_TS(21) or SL6_TS(22) or SL6_TS(23) ;
SL6_row10(49)<=SL6_TS(23) or SL6_TS(24) or SL6_TS(25) ;
SL6_row10(50)<=SL6_TS(25) or SL6_TS(26) or SL6_TS(27) ;
SL6_row10(51)<=SL6_TS(27) or SL6_TS(28) or SL6_TS(29) ;
SL6_row10(52)<=SL6_TS(29) or SL6_TS(30) or SL6_TS(31) ;
SL6_row10(53)<=SL6_TS(31) or SL6_TS(32) or SL6_TS(33) ;
SL6_row10(54)<=SL6_TS(33) or SL6_TS(34) or SL6_TS(35) ;
SL6_row10(55)<=SL6_TS(35) or SL6_TS(36) or SL6_TS(37) ;
SL6_row10(56)<=SL6_TS(37) or SL6_TS(38) or SL6_TS(39) ;
SL6_row10(57)<=SL6_TS(39) or SL6_TS(40) or SL6_TS(41) ;
SL6_row10(58)<=SL6_TS(41) or SL6_TS(42) or SL6_TS(43) ;
SL6_row10(59)<=SL6_TS(43) or SL6_TS(44) or SL6_TS(45) ;
SL6_row10(60)<=SL6_TS(45) or SL6_TS(46) or SL6_TS(47) ;
SL6_row10(61)<=SL6_TS(47) or SL6_TS(48) or SL6_TS(49) ;
SL6_row10(62)<=SL6_TS(49) or SL6_TS(50) or SL6_TS(51) ;
SL6_row10(63)<=SL6_TS(51) or SL6_TS(52) or SL6_TS(53) ;
SL6_row10(64)<=SL6_TS(53) or SL6_TS(54) or SL6_TS(55) ;
SL6_row10(65)<=SL6_TS(55) or SL6_TS(56) or SL6_TS(57) ;
SL6_row10(66)<=SL6_TS(57) or SL6_TS(58) or SL6_TS(59) ;
SL6_row10(67)<=SL6_TS(59) or SL6_TS(60) or SL6_TS(61) ;
SL6_row10(68)<=SL6_TS(61) or SL6_TS(62) or SL6_TS(63) ;
SL6_row10(69)<=SL6_TS(63) or SL6_TS(64) or SL6_TS(65) ;
SL6_row10(70)<=SL6_TS(65) or SL6_TS(66) or SL6_TS(67) ;
SL6_row10(71)<=SL6_TS(67) or SL6_TS(68) or SL6_TS(69) ;
SL6_row10(72)<=SL6_TS(69) or SL6_TS(70) or SL6_TS(71) ;
SL6_row10(73)<=SL6_TS(71) or SL6_TS(72) or SL6_TS(73) ;
SL6_row10(74)<=SL6_TS(73) or SL6_TS(74) or SL6_TS(75) ;
SL6_row10(75)<=SL6_TS(75) or SL6_TS(76) or SL6_TS(77) ;
SL6_row10(76)<=SL6_TS(77) or SL6_TS(78) or SL6_TS(79) ;
SL6_row10(77)<=SL6_TS(79) or SL6_TS(80) or SL6_TS(81) ;
SL6_row10(78)<=SL6_TS(81) or SL6_TS(82) or SL6_TS(83) ;
SL6_row10(79)<=SL6_TS(83) or SL6_TS(84) or SL6_TS(85) ;
SL6_row11(40)<=SL6_TS(4) or SL6_TS(5) or SL6_TS(6) ;
SL6_row11(41)<=SL6_TS(6) or SL6_TS(7) or SL6_TS(8) ;
SL6_row11(42)<=SL6_TS(8) or SL6_TS(9) or SL6_TS(10) ;
SL6_row11(43)<=SL6_TS(10) or SL6_TS(11) or SL6_TS(12) ;
SL6_row11(44)<=SL6_TS(12) or SL6_TS(13) or SL6_TS(14) ;
SL6_row11(45)<=SL6_TS(14) or SL6_TS(15) or SL6_TS(16) ;
SL6_row11(46)<=SL6_TS(16) or SL6_TS(17) or SL6_TS(18) ;
SL6_row11(47)<=SL6_TS(18) or SL6_TS(19) or SL6_TS(20) ;
SL6_row11(48)<=SL6_TS(20) or SL6_TS(21) or SL6_TS(22) ;
SL6_row11(49)<=SL6_TS(22) or SL6_TS(23) or SL6_TS(24) ;
SL6_row11(50)<=SL6_TS(24) or SL6_TS(25) or SL6_TS(26) ;
SL6_row11(51)<=SL6_TS(26) or SL6_TS(27) or SL6_TS(28) ;
SL6_row11(52)<=SL6_TS(28) or SL6_TS(29) or SL6_TS(30) ;
SL6_row11(53)<=SL6_TS(30) or SL6_TS(31) or SL6_TS(32) ;
SL6_row11(54)<=SL6_TS(32) or SL6_TS(33) or SL6_TS(34) ;
SL6_row11(55)<=SL6_TS(34) or SL6_TS(35) or SL6_TS(36) ;
SL6_row11(56)<=SL6_TS(36) or SL6_TS(37) or SL6_TS(38) ;
SL6_row11(57)<=SL6_TS(38) or SL6_TS(39) or SL6_TS(40) ;
SL6_row11(58)<=SL6_TS(40) or SL6_TS(41) or SL6_TS(42) ;
SL6_row11(59)<=SL6_TS(42) or SL6_TS(43) or SL6_TS(44) ;
SL6_row11(60)<=SL6_TS(44) or SL6_TS(45) or SL6_TS(46) ;
SL6_row11(61)<=SL6_TS(46) or SL6_TS(47) or SL6_TS(48) ;
SL6_row11(62)<=SL6_TS(48) or SL6_TS(49) or SL6_TS(50) ;
SL6_row11(63)<=SL6_TS(50) or SL6_TS(51) or SL6_TS(52) ;
SL6_row11(64)<=SL6_TS(52) or SL6_TS(53) or SL6_TS(54) ;
SL6_row11(65)<=SL6_TS(54) or SL6_TS(55) or SL6_TS(56) ;
SL6_row11(66)<=SL6_TS(56) or SL6_TS(57) or SL6_TS(58) ;
SL6_row11(67)<=SL6_TS(58) or SL6_TS(59) or SL6_TS(60) ;
SL6_row11(68)<=SL6_TS(60) or SL6_TS(61) or SL6_TS(62) ;
SL6_row11(69)<=SL6_TS(62) or SL6_TS(63) or SL6_TS(64) ;
SL6_row11(70)<=SL6_TS(64) or SL6_TS(65) or SL6_TS(66) ;
SL6_row11(71)<=SL6_TS(66) or SL6_TS(67) or SL6_TS(68) ;
SL6_row11(72)<=SL6_TS(68) or SL6_TS(69) or SL6_TS(70) ;
SL6_row11(73)<=SL6_TS(70) or SL6_TS(71) or SL6_TS(72) ;
SL6_row11(74)<=SL6_TS(72) or SL6_TS(73) or SL6_TS(74) ;
SL6_row11(75)<=SL6_TS(74) or SL6_TS(75) or SL6_TS(76) ;
SL6_row11(76)<=SL6_TS(76) or SL6_TS(77) or SL6_TS(78) ;
SL6_row11(77)<=SL6_TS(78) or SL6_TS(79) or SL6_TS(80) ;
SL6_row11(78)<=SL6_TS(80) or SL6_TS(81) or SL6_TS(82) ;
SL6_row11(79)<=SL6_TS(82) or SL6_TS(83) or SL6_TS(84) ;
SL6_row12(40)<=SL6_TS(3) or SL6_TS(4) or SL6_TS(5) ;
SL6_row12(41)<=SL6_TS(5) or SL6_TS(6) or SL6_TS(7) ;
SL6_row12(42)<=SL6_TS(7) or SL6_TS(8) or SL6_TS(9) ;
SL6_row12(43)<=SL6_TS(9) or SL6_TS(10) or SL6_TS(11) ;
SL6_row12(44)<=SL6_TS(11) or SL6_TS(12) or SL6_TS(13) ;
SL6_row12(45)<=SL6_TS(13) or SL6_TS(14) or SL6_TS(15) ;
SL6_row12(46)<=SL6_TS(15) or SL6_TS(16) or SL6_TS(17) ;
SL6_row12(47)<=SL6_TS(17) or SL6_TS(18) or SL6_TS(19) ;
SL6_row12(48)<=SL6_TS(19) or SL6_TS(20) or SL6_TS(21) ;
SL6_row12(49)<=SL6_TS(21) or SL6_TS(22) or SL6_TS(23) ;
SL6_row12(50)<=SL6_TS(23) or SL6_TS(24) or SL6_TS(25) ;
SL6_row12(51)<=SL6_TS(25) or SL6_TS(26) or SL6_TS(27) ;
SL6_row12(52)<=SL6_TS(27) or SL6_TS(28) or SL6_TS(29) ;
SL6_row12(53)<=SL6_TS(29) or SL6_TS(30) or SL6_TS(31) ;
SL6_row12(54)<=SL6_TS(31) or SL6_TS(32) or SL6_TS(33) ;
SL6_row12(55)<=SL6_TS(33) or SL6_TS(34) or SL6_TS(35) ;
SL6_row12(56)<=SL6_TS(35) or SL6_TS(36) or SL6_TS(37) ;
SL6_row12(57)<=SL6_TS(37) or SL6_TS(38) or SL6_TS(39) ;
SL6_row12(58)<=SL6_TS(39) or SL6_TS(40) or SL6_TS(41) ;
SL6_row12(59)<=SL6_TS(41) or SL6_TS(42) or SL6_TS(43) ;
SL6_row12(60)<=SL6_TS(43) or SL6_TS(44) or SL6_TS(45) ;
SL6_row12(61)<=SL6_TS(45) or SL6_TS(46) or SL6_TS(47) ;
SL6_row12(62)<=SL6_TS(47) or SL6_TS(48) or SL6_TS(49) ;
SL6_row12(63)<=SL6_TS(49) or SL6_TS(50) or SL6_TS(51) ;
SL6_row12(64)<=SL6_TS(51) or SL6_TS(52) or SL6_TS(53) ;
SL6_row12(65)<=SL6_TS(53) or SL6_TS(54) or SL6_TS(55) ;
SL6_row12(66)<=SL6_TS(55) or SL6_TS(56) or SL6_TS(57) ;
SL6_row12(67)<=SL6_TS(57) or SL6_TS(58) or SL6_TS(59) ;
SL6_row12(68)<=SL6_TS(59) or SL6_TS(60) or SL6_TS(61) ;
SL6_row12(69)<=SL6_TS(61) or SL6_TS(62) or SL6_TS(63) ;
SL6_row12(70)<=SL6_TS(63) or SL6_TS(64) or SL6_TS(65) ;
SL6_row12(71)<=SL6_TS(65) or SL6_TS(66) or SL6_TS(67) ;
SL6_row12(72)<=SL6_TS(67) or SL6_TS(68) or SL6_TS(69) ;
SL6_row12(73)<=SL6_TS(69) or SL6_TS(70) or SL6_TS(71) ;
SL6_row12(74)<=SL6_TS(71) or SL6_TS(72) or SL6_TS(73) ;
SL6_row12(75)<=SL6_TS(73) or SL6_TS(74) or SL6_TS(75) ;
SL6_row12(76)<=SL6_TS(75) or SL6_TS(76) or SL6_TS(77) ;
SL6_row12(77)<=SL6_TS(77) or SL6_TS(78) or SL6_TS(79) ;
SL6_row12(78)<=SL6_TS(79) or SL6_TS(80) or SL6_TS(81) ;
SL6_row12(79)<=SL6_TS(81) or SL6_TS(82) or SL6_TS(83) ;
SL6_row13(40)<=SL6_TS(3) or SL6_TS(4) ;
SL6_row13(41)<=SL6_TS(5) or SL6_TS(6) ;
SL6_row13(42)<=SL6_TS(7) or SL6_TS(8) ;
SL6_row13(43)<=SL6_TS(9) or SL6_TS(10) ;
SL6_row13(44)<=SL6_TS(11) or SL6_TS(12) ;
SL6_row13(45)<=SL6_TS(13) or SL6_TS(14) ;
SL6_row13(46)<=SL6_TS(15) or SL6_TS(16) ;
SL6_row13(47)<=SL6_TS(17) or SL6_TS(18) ;
SL6_row13(48)<=SL6_TS(19) or SL6_TS(20) ;
SL6_row13(49)<=SL6_TS(21) or SL6_TS(22) ;
SL6_row13(50)<=SL6_TS(23) or SL6_TS(24) ;
SL6_row13(51)<=SL6_TS(25) or SL6_TS(26) ;
SL6_row13(52)<=SL6_TS(27) or SL6_TS(28) ;
SL6_row13(53)<=SL6_TS(29) or SL6_TS(30) ;
SL6_row13(54)<=SL6_TS(31) or SL6_TS(32) ;
SL6_row13(55)<=SL6_TS(33) or SL6_TS(34) ;
SL6_row13(56)<=SL6_TS(35) or SL6_TS(36) ;
SL6_row13(57)<=SL6_TS(37) or SL6_TS(38) ;
SL6_row13(58)<=SL6_TS(39) or SL6_TS(40) ;
SL6_row13(59)<=SL6_TS(41) or SL6_TS(42) ;
SL6_row13(60)<=SL6_TS(43) or SL6_TS(44) ;
SL6_row13(61)<=SL6_TS(45) or SL6_TS(46) ;
SL6_row13(62)<=SL6_TS(47) or SL6_TS(48) ;
SL6_row13(63)<=SL6_TS(49) or SL6_TS(50) ;
SL6_row13(64)<=SL6_TS(51) or SL6_TS(52) ;
SL6_row13(65)<=SL6_TS(53) or SL6_TS(54) ;
SL6_row13(66)<=SL6_TS(55) or SL6_TS(56) ;
SL6_row13(67)<=SL6_TS(57) or SL6_TS(58) ;
SL6_row13(68)<=SL6_TS(59) or SL6_TS(60) ;
SL6_row13(69)<=SL6_TS(61) or SL6_TS(62) ;
SL6_row13(70)<=SL6_TS(63) or SL6_TS(64) ;
SL6_row13(71)<=SL6_TS(65) or SL6_TS(66) ;
SL6_row13(72)<=SL6_TS(67) or SL6_TS(68) ;
SL6_row13(73)<=SL6_TS(69) or SL6_TS(70) ;
SL6_row13(74)<=SL6_TS(71) or SL6_TS(72) ;
SL6_row13(75)<=SL6_TS(73) or SL6_TS(74) ;
SL6_row13(76)<=SL6_TS(75) or SL6_TS(76) ;
SL6_row13(77)<=SL6_TS(77) or SL6_TS(78) ;
SL6_row13(78)<=SL6_TS(79) or SL6_TS(80) ;
SL6_row13(79)<=SL6_TS(81) or SL6_TS(82) ;
SL6_row14(40)<=SL6_TS(2) or SL6_TS(3) or SL6_TS(4) ;
SL6_row14(41)<=SL6_TS(4) or SL6_TS(5) or SL6_TS(6) ;
SL6_row14(42)<=SL6_TS(6) or SL6_TS(7) or SL6_TS(8) ;
SL6_row14(43)<=SL6_TS(8) or SL6_TS(9) or SL6_TS(10) ;
SL6_row14(44)<=SL6_TS(10) or SL6_TS(11) or SL6_TS(12) ;
SL6_row14(45)<=SL6_TS(12) or SL6_TS(13) or SL6_TS(14) ;
SL6_row14(46)<=SL6_TS(14) or SL6_TS(15) or SL6_TS(16) ;
SL6_row14(47)<=SL6_TS(16) or SL6_TS(17) or SL6_TS(18) ;
SL6_row14(48)<=SL6_TS(18) or SL6_TS(19) or SL6_TS(20) ;
SL6_row14(49)<=SL6_TS(20) or SL6_TS(21) or SL6_TS(22) ;
SL6_row14(50)<=SL6_TS(22) or SL6_TS(23) or SL6_TS(24) ;
SL6_row14(51)<=SL6_TS(24) or SL6_TS(25) or SL6_TS(26) ;
SL6_row14(52)<=SL6_TS(26) or SL6_TS(27) or SL6_TS(28) ;
SL6_row14(53)<=SL6_TS(28) or SL6_TS(29) or SL6_TS(30) ;
SL6_row14(54)<=SL6_TS(30) or SL6_TS(31) or SL6_TS(32) ;
SL6_row14(55)<=SL6_TS(32) or SL6_TS(33) or SL6_TS(34) ;
SL6_row14(56)<=SL6_TS(34) or SL6_TS(35) or SL6_TS(36) ;
SL6_row14(57)<=SL6_TS(36) or SL6_TS(37) or SL6_TS(38) ;
SL6_row14(58)<=SL6_TS(38) or SL6_TS(39) or SL6_TS(40) ;
SL6_row14(59)<=SL6_TS(40) or SL6_TS(41) or SL6_TS(42) ;
SL6_row14(60)<=SL6_TS(42) or SL6_TS(43) or SL6_TS(44) ;
SL6_row14(61)<=SL6_TS(44) or SL6_TS(45) or SL6_TS(46) ;
SL6_row14(62)<=SL6_TS(46) or SL6_TS(47) or SL6_TS(48) ;
SL6_row14(63)<=SL6_TS(48) or SL6_TS(49) or SL6_TS(50) ;
SL6_row14(64)<=SL6_TS(50) or SL6_TS(51) or SL6_TS(52) ;
SL6_row14(65)<=SL6_TS(52) or SL6_TS(53) or SL6_TS(54) ;
SL6_row14(66)<=SL6_TS(54) or SL6_TS(55) or SL6_TS(56) ;
SL6_row14(67)<=SL6_TS(56) or SL6_TS(57) or SL6_TS(58) ;
SL6_row14(68)<=SL6_TS(58) or SL6_TS(59) or SL6_TS(60) ;
SL6_row14(69)<=SL6_TS(60) or SL6_TS(61) or SL6_TS(62) ;
SL6_row14(70)<=SL6_TS(62) or SL6_TS(63) or SL6_TS(64) ;
SL6_row14(71)<=SL6_TS(64) or SL6_TS(65) or SL6_TS(66) ;
SL6_row14(72)<=SL6_TS(66) or SL6_TS(67) or SL6_TS(68) ;
SL6_row14(73)<=SL6_TS(68) or SL6_TS(69) or SL6_TS(70) ;
SL6_row14(74)<=SL6_TS(70) or SL6_TS(71) or SL6_TS(72) ;
SL6_row14(75)<=SL6_TS(72) or SL6_TS(73) or SL6_TS(74) ;
SL6_row14(76)<=SL6_TS(74) or SL6_TS(75) or SL6_TS(76) ;
SL6_row14(77)<=SL6_TS(76) or SL6_TS(77) or SL6_TS(78) ;
SL6_row14(78)<=SL6_TS(78) or SL6_TS(79) or SL6_TS(80) ;
SL6_row14(79)<=SL6_TS(80) or SL6_TS(81) or SL6_TS(82) ;
SL6_row15(40)<=SL6_TS(2) or SL6_TS(3) ;
SL6_row15(41)<=SL6_TS(4) or SL6_TS(5) ;
SL6_row15(42)<=SL6_TS(6) or SL6_TS(7) ;
SL6_row15(43)<=SL6_TS(8) or SL6_TS(9) ;
SL6_row15(44)<=SL6_TS(10) or SL6_TS(11) ;
SL6_row15(45)<=SL6_TS(12) or SL6_TS(13) ;
SL6_row15(46)<=SL6_TS(14) or SL6_TS(15) ;
SL6_row15(47)<=SL6_TS(16) or SL6_TS(17) ;
SL6_row15(48)<=SL6_TS(18) or SL6_TS(19) ;
SL6_row15(49)<=SL6_TS(20) or SL6_TS(21) ;
SL6_row15(50)<=SL6_TS(22) or SL6_TS(23) ;
SL6_row15(51)<=SL6_TS(24) or SL6_TS(25) ;
SL6_row15(52)<=SL6_TS(26) or SL6_TS(27) ;
SL6_row15(53)<=SL6_TS(28) or SL6_TS(29) ;
SL6_row15(54)<=SL6_TS(30) or SL6_TS(31) ;
SL6_row15(55)<=SL6_TS(32) or SL6_TS(33) ;
SL6_row15(56)<=SL6_TS(34) or SL6_TS(35) ;
SL6_row15(57)<=SL6_TS(36) or SL6_TS(37) ;
SL6_row15(58)<=SL6_TS(38) or SL6_TS(39) ;
SL6_row15(59)<=SL6_TS(40) or SL6_TS(41) ;
SL6_row15(60)<=SL6_TS(42) or SL6_TS(43) ;
SL6_row15(61)<=SL6_TS(44) or SL6_TS(45) ;
SL6_row15(62)<=SL6_TS(46) or SL6_TS(47) ;
SL6_row15(63)<=SL6_TS(48) or SL6_TS(49) ;
SL6_row15(64)<=SL6_TS(50) or SL6_TS(51) ;
SL6_row15(65)<=SL6_TS(52) or SL6_TS(53) ;
SL6_row15(66)<=SL6_TS(54) or SL6_TS(55) ;
SL6_row15(67)<=SL6_TS(56) or SL6_TS(57) ;
SL6_row15(68)<=SL6_TS(58) or SL6_TS(59) ;
SL6_row15(69)<=SL6_TS(60) or SL6_TS(61) ;
SL6_row15(70)<=SL6_TS(62) or SL6_TS(63) ;
SL6_row15(71)<=SL6_TS(64) or SL6_TS(65) ;
SL6_row15(72)<=SL6_TS(66) or SL6_TS(67) ;
SL6_row15(73)<=SL6_TS(68) or SL6_TS(69) ;
SL6_row15(74)<=SL6_TS(70) or SL6_TS(71) ;
SL6_row15(75)<=SL6_TS(72) or SL6_TS(73) ;
SL6_row15(76)<=SL6_TS(74) or SL6_TS(75) ;
SL6_row15(77)<=SL6_TS(76) or SL6_TS(77) ;
SL6_row15(78)<=SL6_TS(78) or SL6_TS(79) ;
SL6_row15(79)<=SL6_TS(80) or SL6_TS(81) ;
SL6_row16(40)<=SL6_TS(2) or SL6_TS(3) ;
SL6_row16(41)<=SL6_TS(4) or SL6_TS(5) ;
SL6_row16(42)<=SL6_TS(6) or SL6_TS(7) ;
SL6_row16(43)<=SL6_TS(8) or SL6_TS(9) ;
SL6_row16(44)<=SL6_TS(10) or SL6_TS(11) ;
SL6_row16(45)<=SL6_TS(12) or SL6_TS(13) ;
SL6_row16(46)<=SL6_TS(14) or SL6_TS(15) ;
SL6_row16(47)<=SL6_TS(16) or SL6_TS(17) ;
SL6_row16(48)<=SL6_TS(18) or SL6_TS(19) ;
SL6_row16(49)<=SL6_TS(20) or SL6_TS(21) ;
SL6_row16(50)<=SL6_TS(22) or SL6_TS(23) ;
SL6_row16(51)<=SL6_TS(24) or SL6_TS(25) ;
SL6_row16(52)<=SL6_TS(26) or SL6_TS(27) ;
SL6_row16(53)<=SL6_TS(28) or SL6_TS(29) ;
SL6_row16(54)<=SL6_TS(30) or SL6_TS(31) ;
SL6_row16(55)<=SL6_TS(32) or SL6_TS(33) ;
SL6_row16(56)<=SL6_TS(34) or SL6_TS(35) ;
SL6_row16(57)<=SL6_TS(36) or SL6_TS(37) ;
SL6_row16(58)<=SL6_TS(38) or SL6_TS(39) ;
SL6_row16(59)<=SL6_TS(40) or SL6_TS(41) ;
SL6_row16(60)<=SL6_TS(42) or SL6_TS(43) ;
SL6_row16(61)<=SL6_TS(44) or SL6_TS(45) ;
SL6_row16(62)<=SL6_TS(46) or SL6_TS(47) ;
SL6_row16(63)<=SL6_TS(48) or SL6_TS(49) ;
SL6_row16(64)<=SL6_TS(50) or SL6_TS(51) ;
SL6_row16(65)<=SL6_TS(52) or SL6_TS(53) ;
SL6_row16(66)<=SL6_TS(54) or SL6_TS(55) ;
SL6_row16(67)<=SL6_TS(56) or SL6_TS(57) ;
SL6_row16(68)<=SL6_TS(58) or SL6_TS(59) ;
SL6_row16(69)<=SL6_TS(60) or SL6_TS(61) ;
SL6_row16(70)<=SL6_TS(62) or SL6_TS(63) ;
SL6_row16(71)<=SL6_TS(64) or SL6_TS(65) ;
SL6_row16(72)<=SL6_TS(66) or SL6_TS(67) ;
SL6_row16(73)<=SL6_TS(68) or SL6_TS(69) ;
SL6_row16(74)<=SL6_TS(70) or SL6_TS(71) ;
SL6_row16(75)<=SL6_TS(72) or SL6_TS(73) ;
SL6_row16(76)<=SL6_TS(74) or SL6_TS(75) ;
SL6_row16(77)<=SL6_TS(76) or SL6_TS(77) ;
SL6_row16(78)<=SL6_TS(78) or SL6_TS(79) ;
SL6_row16(79)<=SL6_TS(80) or SL6_TS(81) ;
 
end Behavioral;

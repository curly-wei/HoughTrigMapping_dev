library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
 
entity UT3_0_SL2_P is
 
Port (
           SL2_row1  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row2  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row3  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row4  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row5  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row6  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row7  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row8  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row9  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row10 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row11 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row12 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row13 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row14 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row15 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_row16 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL2_TS    : in   STD_LOGIC_VECTOR (96 downto 0));
end UT3_0_SL2_P;
 
 
architecture Behavioral of UT3_0_SL2_P is
 
begin
 
SL2_row1(0)<=SL2_TS(39) or SL2_TS(40) or SL2_TS(41) ;
SL2_row1(1)<=SL2_TS(40) or SL2_TS(41) or SL2_TS(42) ;
SL2_row1(2)<=SL2_TS(42) or SL2_TS(43) ;
SL2_row1(3)<=SL2_TS(43) or SL2_TS(44) or SL2_TS(45) ;
SL2_row1(4)<=SL2_TS(44) or SL2_TS(45) or SL2_TS(46) ;
SL2_row1(5)<=SL2_TS(45) or SL2_TS(46) or SL2_TS(47) ;
SL2_row1(6)<=SL2_TS(46) or SL2_TS(47) or SL2_TS(48) ;
SL2_row1(7)<=SL2_TS(48) or SL2_TS(49) ;
SL2_row1(8)<=SL2_TS(49) or SL2_TS(50) or SL2_TS(51) ;
SL2_row1(9)<=SL2_TS(50) or SL2_TS(51) or SL2_TS(52) ;
SL2_row1(10)<=SL2_TS(51) or SL2_TS(52) or SL2_TS(53) ;
SL2_row1(11)<=SL2_TS(52) or SL2_TS(53) or SL2_TS(54) ;
SL2_row1(12)<=SL2_TS(54) or SL2_TS(55) ;
SL2_row1(13)<=SL2_TS(55) or SL2_TS(56) or SL2_TS(57) ;
SL2_row1(14)<=SL2_TS(56) or SL2_TS(57) or SL2_TS(58) ;
SL2_row1(15)<=SL2_TS(57) or SL2_TS(58) or SL2_TS(59) ;
SL2_row1(16)<=SL2_TS(58) or SL2_TS(59) or SL2_TS(60) ;
SL2_row1(17)<=SL2_TS(60) or SL2_TS(61) ;
SL2_row1(18)<=SL2_TS(61) or SL2_TS(62) or SL2_TS(63) ;
SL2_row1(19)<=SL2_TS(62) or SL2_TS(63) or SL2_TS(64) ;
SL2_row1(20)<=SL2_TS(63) or SL2_TS(64) or SL2_TS(65) ;
SL2_row1(21)<=SL2_TS(64) or SL2_TS(65) or SL2_TS(66) ;
SL2_row1(22)<=SL2_TS(66) or SL2_TS(67) ;
SL2_row1(23)<=SL2_TS(67) or SL2_TS(68) or SL2_TS(69) ;
SL2_row1(24)<=SL2_TS(68) or SL2_TS(69) or SL2_TS(70) ;
SL2_row1(25)<=SL2_TS(69) or SL2_TS(70) or SL2_TS(71) ;
SL2_row1(26)<=SL2_TS(70) or SL2_TS(71) or SL2_TS(72) ;
SL2_row1(27)<=SL2_TS(72) or SL2_TS(73) ;
SL2_row1(28)<=SL2_TS(73) or SL2_TS(74) or SL2_TS(75) ;
SL2_row1(29)<=SL2_TS(74) or SL2_TS(75) or SL2_TS(76) ;
SL2_row1(30)<=SL2_TS(75) or SL2_TS(76) or SL2_TS(77) ;
SL2_row1(31)<=SL2_TS(76) or SL2_TS(77) or SL2_TS(78) ;
SL2_row1(32)<=SL2_TS(78) or SL2_TS(79) ;
SL2_row1(33)<=SL2_TS(79) or SL2_TS(80) or SL2_TS(81) ;
SL2_row1(34)<=SL2_TS(80) or SL2_TS(81) or SL2_TS(82) ;
SL2_row1(35)<=SL2_TS(81) or SL2_TS(82) or SL2_TS(83) ;
SL2_row1(36)<=SL2_TS(82) or SL2_TS(83) or SL2_TS(84) ;
SL2_row1(37)<=SL2_TS(84) or SL2_TS(85) ;
SL2_row1(38)<=SL2_TS(85) or SL2_TS(86) or SL2_TS(87) ;
SL2_row1(39)<=SL2_TS(86) or SL2_TS(87) or SL2_TS(88) ;
SL2_row2(0)<=SL2_TS(41) or SL2_TS(42) ;
SL2_row2(1)<=SL2_TS(42) or SL2_TS(43) or SL2_TS(44) ;
SL2_row2(2)<=SL2_TS(43) or SL2_TS(44) or SL2_TS(45) ;
SL2_row2(3)<=SL2_TS(44) or SL2_TS(45) or SL2_TS(46) ;
SL2_row2(4)<=SL2_TS(46) or SL2_TS(47) ;
SL2_row2(5)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row2(6)<=SL2_TS(48) or SL2_TS(49) or SL2_TS(50) ;
SL2_row2(7)<=SL2_TS(49) or SL2_TS(50) or SL2_TS(51) ;
SL2_row2(8)<=SL2_TS(50) or SL2_TS(51) or SL2_TS(52) ;
SL2_row2(9)<=SL2_TS(52) or SL2_TS(53) ;
SL2_row2(10)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row2(11)<=SL2_TS(54) or SL2_TS(55) or SL2_TS(56) ;
SL2_row2(12)<=SL2_TS(55) or SL2_TS(56) or SL2_TS(57) ;
SL2_row2(13)<=SL2_TS(56) or SL2_TS(57) or SL2_TS(58) ;
SL2_row2(14)<=SL2_TS(58) or SL2_TS(59) ;
SL2_row2(15)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row2(16)<=SL2_TS(60) or SL2_TS(61) or SL2_TS(62) ;
SL2_row2(17)<=SL2_TS(61) or SL2_TS(62) or SL2_TS(63) ;
SL2_row2(18)<=SL2_TS(62) or SL2_TS(63) or SL2_TS(64) ;
SL2_row2(19)<=SL2_TS(64) or SL2_TS(65) ;
SL2_row2(20)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row2(21)<=SL2_TS(66) or SL2_TS(67) or SL2_TS(68) ;
SL2_row2(22)<=SL2_TS(67) or SL2_TS(68) or SL2_TS(69) ;
SL2_row2(23)<=SL2_TS(68) or SL2_TS(69) or SL2_TS(70) ;
SL2_row2(24)<=SL2_TS(70) or SL2_TS(71) ;
SL2_row2(25)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row2(26)<=SL2_TS(72) or SL2_TS(73) or SL2_TS(74) ;
SL2_row2(27)<=SL2_TS(73) or SL2_TS(74) or SL2_TS(75) ;
SL2_row2(28)<=SL2_TS(74) or SL2_TS(75) or SL2_TS(76) ;
SL2_row2(29)<=SL2_TS(76) or SL2_TS(77) ;
SL2_row2(30)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row2(31)<=SL2_TS(78) or SL2_TS(79) or SL2_TS(80) ;
SL2_row2(32)<=SL2_TS(79) or SL2_TS(80) or SL2_TS(81) ;
SL2_row2(33)<=SL2_TS(80) or SL2_TS(81) or SL2_TS(82) ;
SL2_row2(34)<=SL2_TS(82) or SL2_TS(83) ;
SL2_row2(35)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row2(36)<=SL2_TS(84) or SL2_TS(85) or SL2_TS(86) ;
SL2_row2(37)<=SL2_TS(85) or SL2_TS(86) or SL2_TS(87) ;
SL2_row2(38)<=SL2_TS(86) or SL2_TS(87) or SL2_TS(88) ;
SL2_row2(39)<=SL2_TS(88) or SL2_TS(89) ;
SL2_row3(0)<=SL2_TS(42) or SL2_TS(43) or SL2_TS(44) ;
SL2_row3(1)<=SL2_TS(43) or SL2_TS(44) or SL2_TS(45) ;
SL2_row3(2)<=SL2_TS(45) or SL2_TS(46) ;
SL2_row3(3)<=SL2_TS(46) or SL2_TS(47) ;
SL2_row3(4)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row3(5)<=SL2_TS(48) or SL2_TS(49) or SL2_TS(50) ;
SL2_row3(6)<=SL2_TS(49) or SL2_TS(50) or SL2_TS(51) ;
SL2_row3(7)<=SL2_TS(51) or SL2_TS(52) ;
SL2_row3(8)<=SL2_TS(52) or SL2_TS(53) ;
SL2_row3(9)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row3(10)<=SL2_TS(54) or SL2_TS(55) or SL2_TS(56) ;
SL2_row3(11)<=SL2_TS(55) or SL2_TS(56) or SL2_TS(57) ;
SL2_row3(12)<=SL2_TS(57) or SL2_TS(58) ;
SL2_row3(13)<=SL2_TS(58) or SL2_TS(59) ;
SL2_row3(14)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row3(15)<=SL2_TS(60) or SL2_TS(61) or SL2_TS(62) ;
SL2_row3(16)<=SL2_TS(61) or SL2_TS(62) or SL2_TS(63) ;
SL2_row3(17)<=SL2_TS(63) or SL2_TS(64) ;
SL2_row3(18)<=SL2_TS(64) or SL2_TS(65) ;
SL2_row3(19)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row3(20)<=SL2_TS(66) or SL2_TS(67) or SL2_TS(68) ;
SL2_row3(21)<=SL2_TS(67) or SL2_TS(68) or SL2_TS(69) ;
SL2_row3(22)<=SL2_TS(69) or SL2_TS(70) ;
SL2_row3(23)<=SL2_TS(70) or SL2_TS(71) ;
SL2_row3(24)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row3(25)<=SL2_TS(72) or SL2_TS(73) or SL2_TS(74) ;
SL2_row3(26)<=SL2_TS(73) or SL2_TS(74) or SL2_TS(75) ;
SL2_row3(27)<=SL2_TS(75) or SL2_TS(76) ;
SL2_row3(28)<=SL2_TS(76) or SL2_TS(77) ;
SL2_row3(29)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row3(30)<=SL2_TS(78) or SL2_TS(79) or SL2_TS(80) ;
SL2_row3(31)<=SL2_TS(79) or SL2_TS(80) or SL2_TS(81) ;
SL2_row3(32)<=SL2_TS(81) or SL2_TS(82) ;
SL2_row3(33)<=SL2_TS(82) or SL2_TS(83) ;
SL2_row3(34)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row3(35)<=SL2_TS(84) or SL2_TS(85) or SL2_TS(86) ;
SL2_row3(36)<=SL2_TS(85) or SL2_TS(86) or SL2_TS(87) ;
SL2_row3(37)<=SL2_TS(87) or SL2_TS(88) ;
SL2_row3(38)<=SL2_TS(88) or SL2_TS(89) ;
SL2_row3(39)<=SL2_TS(89) or SL2_TS(90) ;
SL2_row4(0)<=SL2_TS(43) or SL2_TS(44) or SL2_TS(45) ;
SL2_row4(1)<=SL2_TS(45) or SL2_TS(46) ;
SL2_row4(2)<=SL2_TS(46) or SL2_TS(47) ;
SL2_row4(3)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row4(4)<=SL2_TS(48) or SL2_TS(49) ;
SL2_row4(5)<=SL2_TS(49) or SL2_TS(50) or SL2_TS(51) ;
SL2_row4(6)<=SL2_TS(51) or SL2_TS(52) ;
SL2_row4(7)<=SL2_TS(52) or SL2_TS(53) ;
SL2_row4(8)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row4(9)<=SL2_TS(54) or SL2_TS(55) ;
SL2_row4(10)<=SL2_TS(55) or SL2_TS(56) or SL2_TS(57) ;
SL2_row4(11)<=SL2_TS(57) or SL2_TS(58) ;
SL2_row4(12)<=SL2_TS(58) or SL2_TS(59) ;
SL2_row4(13)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row4(14)<=SL2_TS(60) or SL2_TS(61) ;
SL2_row4(15)<=SL2_TS(61) or SL2_TS(62) or SL2_TS(63) ;
SL2_row4(16)<=SL2_TS(63) or SL2_TS(64) ;
SL2_row4(17)<=SL2_TS(64) or SL2_TS(65) ;
SL2_row4(18)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row4(19)<=SL2_TS(66) or SL2_TS(67) ;
SL2_row4(20)<=SL2_TS(67) or SL2_TS(68) or SL2_TS(69) ;
SL2_row4(21)<=SL2_TS(69) or SL2_TS(70) ;
SL2_row4(22)<=SL2_TS(70) or SL2_TS(71) ;
SL2_row4(23)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row4(24)<=SL2_TS(72) or SL2_TS(73) ;
SL2_row4(25)<=SL2_TS(73) or SL2_TS(74) or SL2_TS(75) ;
SL2_row4(26)<=SL2_TS(75) or SL2_TS(76) ;
SL2_row4(27)<=SL2_TS(76) or SL2_TS(77) ;
SL2_row4(28)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row4(29)<=SL2_TS(78) or SL2_TS(79) ;
SL2_row4(30)<=SL2_TS(79) or SL2_TS(80) or SL2_TS(81) ;
SL2_row4(31)<=SL2_TS(81) or SL2_TS(82) ;
SL2_row4(32)<=SL2_TS(82) or SL2_TS(83) ;
SL2_row4(33)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row4(34)<=SL2_TS(84) or SL2_TS(85) ;
SL2_row4(35)<=SL2_TS(85) or SL2_TS(86) or SL2_TS(87) ;
SL2_row4(36)<=SL2_TS(87) or SL2_TS(88) ;
SL2_row4(37)<=SL2_TS(88) or SL2_TS(89) ;
SL2_row4(38)<=SL2_TS(89) or SL2_TS(90) ;
SL2_row4(39)<=SL2_TS(90) or SL2_TS(91) ;
SL2_row5(0)<=SL2_TS(44) or SL2_TS(45) ;
SL2_row5(1)<=SL2_TS(46) ;
SL2_row5(2)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row5(3)<=SL2_TS(48) or SL2_TS(49) ;
SL2_row5(4)<=SL2_TS(49) or SL2_TS(50) ;
SL2_row5(5)<=SL2_TS(50) or SL2_TS(51) ;
SL2_row5(6)<=SL2_TS(52) ;
SL2_row5(7)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row5(8)<=SL2_TS(54) or SL2_TS(55) ;
SL2_row5(9)<=SL2_TS(55) or SL2_TS(56) ;
SL2_row5(10)<=SL2_TS(56) or SL2_TS(57) ;
SL2_row5(11)<=SL2_TS(58) ;
SL2_row5(12)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row5(13)<=SL2_TS(60) or SL2_TS(61) ;
SL2_row5(14)<=SL2_TS(61) or SL2_TS(62) ;
SL2_row5(15)<=SL2_TS(62) or SL2_TS(63) ;
SL2_row5(16)<=SL2_TS(64) ;
SL2_row5(17)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row5(18)<=SL2_TS(66) or SL2_TS(67) ;
SL2_row5(19)<=SL2_TS(67) or SL2_TS(68) ;
SL2_row5(20)<=SL2_TS(68) or SL2_TS(69) ;
SL2_row5(21)<=SL2_TS(70) ;
SL2_row5(22)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row5(23)<=SL2_TS(72) or SL2_TS(73) ;
SL2_row5(24)<=SL2_TS(73) or SL2_TS(74) ;
SL2_row5(25)<=SL2_TS(74) or SL2_TS(75) ;
SL2_row5(26)<=SL2_TS(76) ;
SL2_row5(27)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row5(28)<=SL2_TS(78) or SL2_TS(79) ;
SL2_row5(29)<=SL2_TS(79) or SL2_TS(80) ;
SL2_row5(30)<=SL2_TS(80) or SL2_TS(81) ;
SL2_row5(31)<=SL2_TS(82) ;
SL2_row5(32)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row5(33)<=SL2_TS(84) or SL2_TS(85) ;
SL2_row5(34)<=SL2_TS(85) or SL2_TS(86) ;
SL2_row5(35)<=SL2_TS(86) or SL2_TS(87) ;
SL2_row5(36)<=SL2_TS(88) ;
SL2_row5(37)<=SL2_TS(89) or SL2_TS(90) ;
SL2_row5(38)<=SL2_TS(90) or SL2_TS(91) ;
SL2_row5(39)<=SL2_TS(91) or SL2_TS(92) ;
SL2_row6(0)<=SL2_TS(45) or SL2_TS(46) ;
SL2_row6(1)<=SL2_TS(46) or SL2_TS(47) ;
SL2_row6(2)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row6(3)<=SL2_TS(49) or SL2_TS(50) ;
SL2_row6(4)<=SL2_TS(50) or SL2_TS(51) ;
SL2_row6(5)<=SL2_TS(51) or SL2_TS(52) ;
SL2_row6(6)<=SL2_TS(52) or SL2_TS(53) ;
SL2_row6(7)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row6(8)<=SL2_TS(55) or SL2_TS(56) ;
SL2_row6(9)<=SL2_TS(56) or SL2_TS(57) ;
SL2_row6(10)<=SL2_TS(57) or SL2_TS(58) ;
SL2_row6(11)<=SL2_TS(58) or SL2_TS(59) ;
SL2_row6(12)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row6(13)<=SL2_TS(61) or SL2_TS(62) ;
SL2_row6(14)<=SL2_TS(62) or SL2_TS(63) ;
SL2_row6(15)<=SL2_TS(63) or SL2_TS(64) ;
SL2_row6(16)<=SL2_TS(64) or SL2_TS(65) ;
SL2_row6(17)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row6(18)<=SL2_TS(67) or SL2_TS(68) ;
SL2_row6(19)<=SL2_TS(68) or SL2_TS(69) ;
SL2_row6(20)<=SL2_TS(69) or SL2_TS(70) ;
SL2_row6(21)<=SL2_TS(70) or SL2_TS(71) ;
SL2_row6(22)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row6(23)<=SL2_TS(73) or SL2_TS(74) ;
SL2_row6(24)<=SL2_TS(74) or SL2_TS(75) ;
SL2_row6(25)<=SL2_TS(75) or SL2_TS(76) ;
SL2_row6(26)<=SL2_TS(76) or SL2_TS(77) ;
SL2_row6(27)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row6(28)<=SL2_TS(79) or SL2_TS(80) ;
SL2_row6(29)<=SL2_TS(80) or SL2_TS(81) ;
SL2_row6(30)<=SL2_TS(81) or SL2_TS(82) ;
SL2_row6(31)<=SL2_TS(82) or SL2_TS(83) ;
SL2_row6(32)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row6(33)<=SL2_TS(85) or SL2_TS(86) ;
SL2_row6(34)<=SL2_TS(86) or SL2_TS(87) ;
SL2_row6(35)<=SL2_TS(87) or SL2_TS(88) ;
SL2_row6(36)<=SL2_TS(88) or SL2_TS(89) ;
SL2_row6(37)<=SL2_TS(89) or SL2_TS(90) ;
SL2_row6(38)<=SL2_TS(91) or SL2_TS(92) ;
SL2_row6(39)<=SL2_TS(92) or SL2_TS(93) ;
SL2_row7(0)<=SL2_TS(46) ;
SL2_row7(1)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row7(2)<=SL2_TS(48) or SL2_TS(49) ;
SL2_row7(3)<=SL2_TS(49) or SL2_TS(50) ;
SL2_row7(4)<=SL2_TS(51) ;
SL2_row7(5)<=SL2_TS(52) ;
SL2_row7(6)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row7(7)<=SL2_TS(54) or SL2_TS(55) ;
SL2_row7(8)<=SL2_TS(55) or SL2_TS(56) ;
SL2_row7(9)<=SL2_TS(57) ;
SL2_row7(10)<=SL2_TS(58) ;
SL2_row7(11)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row7(12)<=SL2_TS(60) or SL2_TS(61) ;
SL2_row7(13)<=SL2_TS(61) or SL2_TS(62) ;
SL2_row7(14)<=SL2_TS(63) ;
SL2_row7(15)<=SL2_TS(64) ;
SL2_row7(16)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row7(17)<=SL2_TS(66) or SL2_TS(67) ;
SL2_row7(18)<=SL2_TS(67) or SL2_TS(68) ;
SL2_row7(19)<=SL2_TS(69) ;
SL2_row7(20)<=SL2_TS(70) ;
SL2_row7(21)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row7(22)<=SL2_TS(72) or SL2_TS(73) ;
SL2_row7(23)<=SL2_TS(73) or SL2_TS(74) ;
SL2_row7(24)<=SL2_TS(75) ;
SL2_row7(25)<=SL2_TS(76) ;
SL2_row7(26)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row7(27)<=SL2_TS(78) or SL2_TS(79) ;
SL2_row7(28)<=SL2_TS(79) or SL2_TS(80) ;
SL2_row7(29)<=SL2_TS(81) ;
SL2_row7(30)<=SL2_TS(82) ;
SL2_row7(31)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row7(32)<=SL2_TS(84) or SL2_TS(85) ;
SL2_row7(33)<=SL2_TS(85) or SL2_TS(86) ;
SL2_row7(34)<=SL2_TS(87) ;
SL2_row7(35)<=SL2_TS(88) ;
SL2_row7(36)<=SL2_TS(89) or SL2_TS(90) ;
SL2_row7(37)<=SL2_TS(90) or SL2_TS(91) ;
SL2_row7(38)<=SL2_TS(91) or SL2_TS(92) ;
SL2_row7(39)<=SL2_TS(93) ;
SL2_row8(0)<=SL2_TS(46) or SL2_TS(47) ;
SL2_row8(1)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row8(2)<=SL2_TS(49) ;
SL2_row8(3)<=SL2_TS(50) ;
SL2_row8(4)<=SL2_TS(51) or SL2_TS(52) ;
SL2_row8(5)<=SL2_TS(52) or SL2_TS(53) ;
SL2_row8(6)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row8(7)<=SL2_TS(55) ;
SL2_row8(8)<=SL2_TS(56) ;
SL2_row8(9)<=SL2_TS(57) or SL2_TS(58) ;
SL2_row8(10)<=SL2_TS(58) or SL2_TS(59) ;
SL2_row8(11)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row8(12)<=SL2_TS(61) ;
SL2_row8(13)<=SL2_TS(62) ;
SL2_row8(14)<=SL2_TS(63) or SL2_TS(64) ;
SL2_row8(15)<=SL2_TS(64) or SL2_TS(65) ;
SL2_row8(16)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row8(17)<=SL2_TS(67) ;
SL2_row8(18)<=SL2_TS(68) ;
SL2_row8(19)<=SL2_TS(69) or SL2_TS(70) ;
SL2_row8(20)<=SL2_TS(70) or SL2_TS(71) ;
SL2_row8(21)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row8(22)<=SL2_TS(73) ;
SL2_row8(23)<=SL2_TS(74) ;
SL2_row8(24)<=SL2_TS(75) or SL2_TS(76) ;
SL2_row8(25)<=SL2_TS(76) or SL2_TS(77) ;
SL2_row8(26)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row8(27)<=SL2_TS(79) ;
SL2_row8(28)<=SL2_TS(80) ;
SL2_row8(29)<=SL2_TS(81) or SL2_TS(82) ;
SL2_row8(30)<=SL2_TS(82) or SL2_TS(83) ;
SL2_row8(31)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row8(32)<=SL2_TS(85) ;
SL2_row8(33)<=SL2_TS(86) ;
SL2_row8(34)<=SL2_TS(87) or SL2_TS(88) ;
SL2_row8(35)<=SL2_TS(88) or SL2_TS(89) ;
SL2_row8(36)<=SL2_TS(89) or SL2_TS(90) ;
SL2_row8(37)<=SL2_TS(91) ;
SL2_row8(38)<=SL2_TS(92) ;
SL2_row8(39)<=SL2_TS(93) or SL2_TS(94) ;
SL2_row9(0)<=SL2_TS(47) ;
SL2_row9(1)<=SL2_TS(48) ;
SL2_row9(2)<=SL2_TS(49) or SL2_TS(50) ;
SL2_row9(3)<=SL2_TS(50) or SL2_TS(51) ;
SL2_row9(4)<=SL2_TS(51) or SL2_TS(52) ;
SL2_row9(5)<=SL2_TS(53) ;
SL2_row9(6)<=SL2_TS(54) ;
SL2_row9(7)<=SL2_TS(55) or SL2_TS(56) ;
SL2_row9(8)<=SL2_TS(56) or SL2_TS(57) ;
SL2_row9(9)<=SL2_TS(57) or SL2_TS(58) ;
SL2_row9(10)<=SL2_TS(59) ;
SL2_row9(11)<=SL2_TS(60) ;
SL2_row9(12)<=SL2_TS(61) or SL2_TS(62) ;
SL2_row9(13)<=SL2_TS(62) or SL2_TS(63) ;
SL2_row9(14)<=SL2_TS(63) or SL2_TS(64) ;
SL2_row9(15)<=SL2_TS(65) ;
SL2_row9(16)<=SL2_TS(66) ;
SL2_row9(17)<=SL2_TS(67) or SL2_TS(68) ;
SL2_row9(18)<=SL2_TS(68) or SL2_TS(69) ;
SL2_row9(19)<=SL2_TS(69) or SL2_TS(70) ;
SL2_row9(20)<=SL2_TS(71) ;
SL2_row9(21)<=SL2_TS(72) ;
SL2_row9(22)<=SL2_TS(73) or SL2_TS(74) ;
SL2_row9(23)<=SL2_TS(74) or SL2_TS(75) ;
SL2_row9(24)<=SL2_TS(75) or SL2_TS(76) ;
SL2_row9(25)<=SL2_TS(77) ;
SL2_row9(26)<=SL2_TS(78) ;
SL2_row9(27)<=SL2_TS(79) or SL2_TS(80) ;
SL2_row9(28)<=SL2_TS(80) or SL2_TS(81) ;
SL2_row9(29)<=SL2_TS(81) or SL2_TS(82) ;
SL2_row9(30)<=SL2_TS(83) ;
SL2_row9(31)<=SL2_TS(84) ;
SL2_row9(32)<=SL2_TS(85) or SL2_TS(86) ;
SL2_row9(33)<=SL2_TS(86) or SL2_TS(87) ;
SL2_row9(34)<=SL2_TS(87) or SL2_TS(88) ;
SL2_row9(35)<=SL2_TS(89) ;
SL2_row9(36)<=SL2_TS(90) ;
SL2_row9(37)<=SL2_TS(91) or SL2_TS(92) ;
SL2_row9(38)<=SL2_TS(92) or SL2_TS(93) ;
SL2_row9(39)<=SL2_TS(93) or SL2_TS(94) ;
SL2_row10(0)<=SL2_TS(47) ;
SL2_row10(1)<=SL2_TS(48) or SL2_TS(49) ;
SL2_row10(2)<=SL2_TS(49) or SL2_TS(50) ;
SL2_row10(3)<=SL2_TS(51) ;
SL2_row10(4)<=SL2_TS(52) ;
SL2_row10(5)<=SL2_TS(53) ;
SL2_row10(6)<=SL2_TS(54) or SL2_TS(55) ;
SL2_row10(7)<=SL2_TS(55) or SL2_TS(56) ;
SL2_row10(8)<=SL2_TS(57) ;
SL2_row10(9)<=SL2_TS(58) ;
SL2_row10(10)<=SL2_TS(59) ;
SL2_row10(11)<=SL2_TS(60) or SL2_TS(61) ;
SL2_row10(12)<=SL2_TS(61) or SL2_TS(62) ;
SL2_row10(13)<=SL2_TS(63) ;
SL2_row10(14)<=SL2_TS(64) ;
SL2_row10(15)<=SL2_TS(65) ;
SL2_row10(16)<=SL2_TS(66) or SL2_TS(67) ;
SL2_row10(17)<=SL2_TS(67) or SL2_TS(68) ;
SL2_row10(18)<=SL2_TS(69) ;
SL2_row10(19)<=SL2_TS(70) ;
SL2_row10(20)<=SL2_TS(71) ;
SL2_row10(21)<=SL2_TS(72) or SL2_TS(73) ;
SL2_row10(22)<=SL2_TS(73) or SL2_TS(74) ;
SL2_row10(23)<=SL2_TS(75) ;
SL2_row10(24)<=SL2_TS(76) ;
SL2_row10(25)<=SL2_TS(77) ;
SL2_row10(26)<=SL2_TS(78) or SL2_TS(79) ;
SL2_row10(27)<=SL2_TS(79) or SL2_TS(80) ;
SL2_row10(28)<=SL2_TS(81) ;
SL2_row10(29)<=SL2_TS(82) ;
SL2_row10(30)<=SL2_TS(83) ;
SL2_row10(31)<=SL2_TS(84) or SL2_TS(85) ;
SL2_row10(32)<=SL2_TS(85) or SL2_TS(86) ;
SL2_row10(33)<=SL2_TS(87) ;
SL2_row10(34)<=SL2_TS(88) ;
SL2_row10(35)<=SL2_TS(89) ;
SL2_row10(36)<=SL2_TS(90) or SL2_TS(91) ;
SL2_row10(37)<=SL2_TS(91) or SL2_TS(92) ;
SL2_row10(38)<=SL2_TS(93) ;
SL2_row10(39)<=SL2_TS(94) ;
SL2_row11(0)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row11(1)<=SL2_TS(48) or SL2_TS(49) ;
SL2_row11(2)<=SL2_TS(50) ;
SL2_row11(3)<=SL2_TS(51) ;
SL2_row11(4)<=SL2_TS(52) ;
SL2_row11(5)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row11(6)<=SL2_TS(54) or SL2_TS(55) ;
SL2_row11(7)<=SL2_TS(56) ;
SL2_row11(8)<=SL2_TS(57) ;
SL2_row11(9)<=SL2_TS(58) ;
SL2_row11(10)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row11(11)<=SL2_TS(60) or SL2_TS(61) ;
SL2_row11(12)<=SL2_TS(62) ;
SL2_row11(13)<=SL2_TS(63) ;
SL2_row11(14)<=SL2_TS(64) ;
SL2_row11(15)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row11(16)<=SL2_TS(66) or SL2_TS(67) ;
SL2_row11(17)<=SL2_TS(68) ;
SL2_row11(18)<=SL2_TS(69) ;
SL2_row11(19)<=SL2_TS(70) ;
SL2_row11(20)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row11(21)<=SL2_TS(72) or SL2_TS(73) ;
SL2_row11(22)<=SL2_TS(74) ;
SL2_row11(23)<=SL2_TS(75) ;
SL2_row11(24)<=SL2_TS(76) ;
SL2_row11(25)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row11(26)<=SL2_TS(78) or SL2_TS(79) ;
SL2_row11(27)<=SL2_TS(80) ;
SL2_row11(28)<=SL2_TS(81) ;
SL2_row11(29)<=SL2_TS(82) ;
SL2_row11(30)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row11(31)<=SL2_TS(84) or SL2_TS(85) ;
SL2_row11(32)<=SL2_TS(86) ;
SL2_row11(33)<=SL2_TS(87) ;
SL2_row11(34)<=SL2_TS(88) ;
SL2_row11(35)<=SL2_TS(89) or SL2_TS(90) ;
SL2_row11(36)<=SL2_TS(90) or SL2_TS(91) ;
SL2_row11(37)<=SL2_TS(92) ;
SL2_row11(38)<=SL2_TS(93) ;
SL2_row11(39)<=SL2_TS(94) ;
SL2_row12(0)<=SL2_TS(47) or SL2_TS(48) ;
SL2_row12(1)<=SL2_TS(49) ;
SL2_row12(2)<=SL2_TS(50) ;
SL2_row12(3)<=SL2_TS(51) ;
SL2_row12(4)<=SL2_TS(52) or SL2_TS(53) ;
SL2_row12(5)<=SL2_TS(53) or SL2_TS(54) ;
SL2_row12(6)<=SL2_TS(55) ;
SL2_row12(7)<=SL2_TS(56) ;
SL2_row12(8)<=SL2_TS(57) ;
SL2_row12(9)<=SL2_TS(58) or SL2_TS(59) ;
SL2_row12(10)<=SL2_TS(59) or SL2_TS(60) ;
SL2_row12(11)<=SL2_TS(61) ;
SL2_row12(12)<=SL2_TS(62) ;
SL2_row12(13)<=SL2_TS(63) ;
SL2_row12(14)<=SL2_TS(64) or SL2_TS(65) ;
SL2_row12(15)<=SL2_TS(65) or SL2_TS(66) ;
SL2_row12(16)<=SL2_TS(67) ;
SL2_row12(17)<=SL2_TS(68) ;
SL2_row12(18)<=SL2_TS(69) ;
SL2_row12(19)<=SL2_TS(70) or SL2_TS(71) ;
SL2_row12(20)<=SL2_TS(71) or SL2_TS(72) ;
SL2_row12(21)<=SL2_TS(73) ;
SL2_row12(22)<=SL2_TS(74) ;
SL2_row12(23)<=SL2_TS(75) ;
SL2_row12(24)<=SL2_TS(76) or SL2_TS(77) ;
SL2_row12(25)<=SL2_TS(77) or SL2_TS(78) ;
SL2_row12(26)<=SL2_TS(79) ;
SL2_row12(27)<=SL2_TS(80) ;
SL2_row12(28)<=SL2_TS(81) ;
SL2_row12(29)<=SL2_TS(82) or SL2_TS(83) ;
SL2_row12(30)<=SL2_TS(83) or SL2_TS(84) ;
SL2_row12(31)<=SL2_TS(85) ;
SL2_row12(32)<=SL2_TS(86) ;
SL2_row12(33)<=SL2_TS(87) ;
SL2_row12(34)<=SL2_TS(88) or SL2_TS(89) ;
SL2_row12(35)<=SL2_TS(89) or SL2_TS(90) ;
SL2_row12(36)<=SL2_TS(91) ;
SL2_row12(37)<=SL2_TS(92) ;
SL2_row12(38)<=SL2_TS(93) ;
SL2_row12(39)<=SL2_TS(94) or SL2_TS(95) ;
SL2_row13(0)<=SL2_TS(48) ;
SL2_row13(1)<=SL2_TS(49) ;
SL2_row13(2)<=SL2_TS(50) ;
SL2_row13(3)<=SL2_TS(51) or SL2_TS(52) ;
SL2_row13(4)<=SL2_TS(52) or SL2_TS(53) ;
SL2_row13(5)<=SL2_TS(54) ;
SL2_row13(6)<=SL2_TS(55) ;
SL2_row13(7)<=SL2_TS(56) ;
SL2_row13(8)<=SL2_TS(57) or SL2_TS(58) ;
SL2_row13(9)<=SL2_TS(58) or SL2_TS(59) ;
SL2_row13(10)<=SL2_TS(60) ;
SL2_row13(11)<=SL2_TS(61) ;
SL2_row13(12)<=SL2_TS(62) ;
SL2_row13(13)<=SL2_TS(63) or SL2_TS(64) ;
SL2_row13(14)<=SL2_TS(64) or SL2_TS(65) ;
SL2_row13(15)<=SL2_TS(66) ;
SL2_row13(16)<=SL2_TS(67) ;
SL2_row13(17)<=SL2_TS(68) ;
SL2_row13(18)<=SL2_TS(69) or SL2_TS(70) ;
SL2_row13(19)<=SL2_TS(70) or SL2_TS(71) ;
SL2_row13(20)<=SL2_TS(72) ;
SL2_row13(21)<=SL2_TS(73) ;
SL2_row13(22)<=SL2_TS(74) ;
SL2_row13(23)<=SL2_TS(75) or SL2_TS(76) ;
SL2_row13(24)<=SL2_TS(76) or SL2_TS(77) ;
SL2_row13(25)<=SL2_TS(78) ;
SL2_row13(26)<=SL2_TS(79) ;
SL2_row13(27)<=SL2_TS(80) ;
SL2_row13(28)<=SL2_TS(81) or SL2_TS(82) ;
SL2_row13(29)<=SL2_TS(82) or SL2_TS(83) ;
SL2_row13(30)<=SL2_TS(84) ;
SL2_row13(31)<=SL2_TS(85) ;
SL2_row13(32)<=SL2_TS(86) ;
SL2_row13(33)<=SL2_TS(87) or SL2_TS(88) ;
SL2_row13(34)<=SL2_TS(88) or SL2_TS(89) ;
SL2_row13(35)<=SL2_TS(90) ;
SL2_row13(36)<=SL2_TS(91) ;
SL2_row13(37)<=SL2_TS(92) ;
SL2_row13(38)<=SL2_TS(93) or SL2_TS(94) ;
SL2_row13(39)<=SL2_TS(94) or SL2_TS(95) ;
SL2_row14(0)<=SL2_TS(48) ;
SL2_row14(1)<=SL2_TS(49) ;
SL2_row14(2)<=SL2_TS(50) or SL2_TS(51) ;
SL2_row14(3)<=SL2_TS(51) or SL2_TS(52) ;
SL2_row14(4)<=SL2_TS(53) ;
SL2_row14(5)<=SL2_TS(54) ;
SL2_row14(6)<=SL2_TS(55) ;
SL2_row14(7)<=SL2_TS(56) or SL2_TS(57) ;
SL2_row14(8)<=SL2_TS(57) or SL2_TS(58) ;
SL2_row14(9)<=SL2_TS(59) ;
SL2_row14(10)<=SL2_TS(60) ;
SL2_row14(11)<=SL2_TS(61) ;
SL2_row14(12)<=SL2_TS(62) or SL2_TS(63) ;
SL2_row14(13)<=SL2_TS(63) or SL2_TS(64) ;
SL2_row14(14)<=SL2_TS(65) ;
SL2_row14(15)<=SL2_TS(66) ;
SL2_row14(16)<=SL2_TS(67) ;
SL2_row14(17)<=SL2_TS(68) or SL2_TS(69) ;
SL2_row14(18)<=SL2_TS(69) or SL2_TS(70) ;
SL2_row14(19)<=SL2_TS(71) ;
SL2_row14(20)<=SL2_TS(72) ;
SL2_row14(21)<=SL2_TS(73) ;
SL2_row14(22)<=SL2_TS(74) or SL2_TS(75) ;
SL2_row14(23)<=SL2_TS(75) or SL2_TS(76) ;
SL2_row14(24)<=SL2_TS(77) ;
SL2_row14(25)<=SL2_TS(78) ;
SL2_row14(26)<=SL2_TS(79) ;
SL2_row14(27)<=SL2_TS(80) or SL2_TS(81) ;
SL2_row14(28)<=SL2_TS(81) or SL2_TS(82) ;
SL2_row14(29)<=SL2_TS(83) ;
SL2_row14(30)<=SL2_TS(84) ;
SL2_row14(31)<=SL2_TS(85) ;
SL2_row14(32)<=SL2_TS(86) or SL2_TS(87) ;
SL2_row14(33)<=SL2_TS(87) or SL2_TS(88) ;
SL2_row14(34)<=SL2_TS(89) ;
SL2_row14(35)<=SL2_TS(90) ;
SL2_row14(36)<=SL2_TS(91) ;
SL2_row14(37)<=SL2_TS(92) or SL2_TS(93) ;
SL2_row14(38)<=SL2_TS(93) or SL2_TS(94) ;
SL2_row14(39)<=SL2_TS(95) ;
SL2_row15(0)<=SL2_TS(48) ;
SL2_row15(1)<=SL2_TS(49) ;
SL2_row15(2)<=SL2_TS(50) or SL2_TS(51) ;
SL2_row15(3)<=SL2_TS(52) ;
SL2_row15(4)<=SL2_TS(53) ;
SL2_row15(5)<=SL2_TS(54) ;
SL2_row15(6)<=SL2_TS(55) ;
SL2_row15(7)<=SL2_TS(56) or SL2_TS(57) ;
SL2_row15(8)<=SL2_TS(58) ;
SL2_row15(9)<=SL2_TS(59) ;
SL2_row15(10)<=SL2_TS(60) ;
SL2_row15(11)<=SL2_TS(61) ;
SL2_row15(12)<=SL2_TS(62) or SL2_TS(63) ;
SL2_row15(13)<=SL2_TS(64) ;
SL2_row15(14)<=SL2_TS(65) ;
SL2_row15(15)<=SL2_TS(66) ;
SL2_row15(16)<=SL2_TS(67) ;
SL2_row15(17)<=SL2_TS(68) or SL2_TS(69) ;
SL2_row15(18)<=SL2_TS(70) ;
SL2_row15(19)<=SL2_TS(71) ;
SL2_row15(20)<=SL2_TS(72) ;
SL2_row15(21)<=SL2_TS(73) ;
SL2_row15(22)<=SL2_TS(74) or SL2_TS(75) ;
SL2_row15(23)<=SL2_TS(76) ;
SL2_row15(24)<=SL2_TS(77) ;
SL2_row15(25)<=SL2_TS(78) ;
SL2_row15(26)<=SL2_TS(79) ;
SL2_row15(27)<=SL2_TS(80) or SL2_TS(81) ;
SL2_row15(28)<=SL2_TS(82) ;
SL2_row15(29)<=SL2_TS(83) ;
SL2_row15(30)<=SL2_TS(84) ;
SL2_row15(31)<=SL2_TS(85) ;
SL2_row15(32)<=SL2_TS(86) or SL2_TS(87) ;
SL2_row15(33)<=SL2_TS(88) ;
SL2_row15(34)<=SL2_TS(89) ;
SL2_row15(35)<=SL2_TS(90) ;
SL2_row15(36)<=SL2_TS(91) ;
SL2_row15(37)<=SL2_TS(92) or SL2_TS(93) ;
SL2_row15(38)<=SL2_TS(94) ;
SL2_row15(39)<=SL2_TS(95) ;
SL2_row16(0)<=SL2_TS(48) ;
SL2_row16(1)<=SL2_TS(49) or SL2_TS(50) ;
SL2_row16(2)<=SL2_TS(50) or SL2_TS(51) ;
SL2_row16(3)<=SL2_TS(52) ;
SL2_row16(4)<=SL2_TS(53) ;
SL2_row16(5)<=SL2_TS(54) ;
SL2_row16(6)<=SL2_TS(55) or SL2_TS(56) ;
SL2_row16(7)<=SL2_TS(56) or SL2_TS(57) ;
SL2_row16(8)<=SL2_TS(58) ;
SL2_row16(9)<=SL2_TS(59) ;
SL2_row16(10)<=SL2_TS(60) ;
SL2_row16(11)<=SL2_TS(61) or SL2_TS(62) ;
SL2_row16(12)<=SL2_TS(62) or SL2_TS(63) ;
SL2_row16(13)<=SL2_TS(64) ;
SL2_row16(14)<=SL2_TS(65) ;
SL2_row16(15)<=SL2_TS(66) ;
SL2_row16(16)<=SL2_TS(67) or SL2_TS(68) ;
SL2_row16(17)<=SL2_TS(68) or SL2_TS(69) ;
SL2_row16(18)<=SL2_TS(70) ;
SL2_row16(19)<=SL2_TS(71) ;
SL2_row16(20)<=SL2_TS(72) ;
SL2_row16(21)<=SL2_TS(73) or SL2_TS(74) ;
SL2_row16(22)<=SL2_TS(74) or SL2_TS(75) ;
SL2_row16(23)<=SL2_TS(76) ;
SL2_row16(24)<=SL2_TS(77) ;
SL2_row16(25)<=SL2_TS(78) ;
SL2_row16(26)<=SL2_TS(79) or SL2_TS(80) ;
SL2_row16(27)<=SL2_TS(80) or SL2_TS(81) ;
SL2_row16(28)<=SL2_TS(82) ;
SL2_row16(29)<=SL2_TS(83) ;
SL2_row16(30)<=SL2_TS(84) ;
SL2_row16(31)<=SL2_TS(85) or SL2_TS(86) ;
SL2_row16(32)<=SL2_TS(86) or SL2_TS(87) ;
SL2_row16(33)<=SL2_TS(88) ;
SL2_row16(34)<=SL2_TS(89) ;
SL2_row16(35)<=SL2_TS(90) ;
SL2_row16(36)<=SL2_TS(91) or SL2_TS(92) ;
SL2_row16(37)<=SL2_TS(92) or SL2_TS(93) ;
SL2_row16(38)<=SL2_TS(94) ;
SL2_row16(39)<=SL2_TS(95) ;
 
end Behavioral;

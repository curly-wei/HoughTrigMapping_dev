library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
 
entity UT3_0_SL0 is
 
Port (
           SL0_map : out SL_map;
           SL0_TS  : in  SL_HIT (NumTSF0 downto 0)
           );
end UT3_0_SL0;
 
 
architecture Behavioral of UT3_0_SL0 is
 
begin
 
SL0_map(0)(0) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(0)(1) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(0)(2) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(0)(3) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(0)(4) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(0)(5) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(0)(6) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(0)(7) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(0)(8) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(0)(9) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(0)(10) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(0)(11) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(0)(12) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(0)(13) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(0)(14) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(0)(15) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(0)(16) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(0)(17) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(0)(18) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(0)(19) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(0)(20) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(0)(21) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(0)(22) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(0)(23) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(0)(24) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(0)(25) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(0)(26) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(0)(27) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(0)(28) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(0)(29) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(0)(30) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(0)(31) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(0)(32) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(0)(33) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(0)(34) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(0)(35) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(0)(36) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(0)(37) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(0)(38) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(0)(39) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(0)(40) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(0)(41) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(0)(42) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(0)(43) <= SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1);
SL0_map(0)(44) <= SL0_TSHit(66)(3) or SL0_TSHit(66)(2) or SL0_TSHit(67)(1);
SL0_map(0)(45) <= SL0_TSHit(67)(3) or SL0_TSHit(67)(2) or SL0_TSHit(68)(1);
SL0_map(1)(0) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(1)(1) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(1)(2) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(1)(3) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(1)(4) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(1)(5) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(1)(6) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(1)(7) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(1)(8) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(1)(9) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(1)(10) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(1)(11) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(1)(12) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(1)(13) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(1)(14) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(1)(15) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(1)(16) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(1)(17) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(1)(18) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(1)(19) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(1)(20) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(1)(21) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(1)(22) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(1)(23) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(1)(24) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(1)(25) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(1)(26) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(1)(27) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(1)(28) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(1)(29) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(1)(30) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(1)(31) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(1)(32) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(1)(33) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(1)(34) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(1)(35) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(1)(36) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(1)(37) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(1)(38) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(1)(39) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(1)(40) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(1)(41) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(1)(42) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(1)(43) <= SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1);
SL0_map(1)(44) <= SL0_TSHit(66)(3) or SL0_TSHit(66)(2) or SL0_TSHit(67)(1);
SL0_map(1)(45) <= SL0_TSHit(67)(3) or SL0_TSHit(67)(2) or SL0_TSHit(68)(1);
SL0_map(2)(0) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(2)(1) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(2)(2) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(2)(3) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(2)(4) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(2)(5) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(2)(6) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(2)(7) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(2)(8) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(2)(9) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(2)(10) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(2)(11) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(2)(12) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(2)(13) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(2)(14) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(2)(15) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(2)(16) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(2)(17) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(2)(18) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(2)(19) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(2)(20) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(2)(21) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(2)(22) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(2)(23) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(2)(24) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(2)(25) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(2)(26) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(2)(27) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(2)(28) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(2)(29) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(2)(30) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(2)(31) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(2)(32) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(2)(33) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(2)(34) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(2)(35) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(2)(36) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(2)(37) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(2)(38) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(2)(39) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(2)(40) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(2)(41) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(2)(42) <= SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(2)(43) <= SL0_TSHit(64)(2) or SL0_TSHit(65)(1) or SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1);
SL0_map(2)(44) <= SL0_TSHit(65)(2) or SL0_TSHit(66)(1) or SL0_TSHit(66)(3) or SL0_TSHit(66)(2) or SL0_TSHit(67)(1);
SL0_map(2)(45) <= SL0_TSHit(66)(2) or SL0_TSHit(67)(1) or SL0_TSHit(67)(3) or SL0_TSHit(67)(2) or SL0_TSHit(68)(1);
SL0_map(3)(0) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(3)(1) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(3)(2) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(3)(3) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(3)(4) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(3)(5) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(3)(6) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(3)(7) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(3)(8) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(3)(9) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(3)(10) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(3)(11) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(3)(12) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(3)(13) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(3)(14) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(3)(15) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(3)(16) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(3)(17) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(3)(18) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(3)(19) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(3)(20) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(3)(21) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(3)(22) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(3)(23) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(3)(24) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(3)(25) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(3)(26) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(3)(27) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(3)(28) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(3)(29) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(3)(30) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(3)(31) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(3)(32) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(3)(33) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(3)(34) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(3)(35) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(3)(36) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(3)(37) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(3)(38) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(3)(39) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(3)(40) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(3)(41) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(3)(42) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3);
SL0_map(3)(43) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1) or SL0_TSHit(65)(3);
SL0_map(3)(44) <= SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1) or SL0_TSHit(66)(3);
SL0_map(3)(45) <= SL0_TSHit(66)(3) or SL0_TSHit(66)(2) or SL0_TSHit(67)(1) or SL0_TSHit(67)(3);
SL0_map(4)(0) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(4)(1) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(4)(2) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(4)(3) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(4)(4) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(4)(5) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(4)(6) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(4)(7) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(4)(8) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(4)(9) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(4)(10) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(4)(11) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(4)(12) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(4)(13) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(4)(14) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(4)(15) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(4)(16) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(4)(17) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(4)(18) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(4)(19) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(4)(20) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(4)(21) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(4)(22) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(4)(23) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(4)(24) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(4)(25) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(4)(26) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(4)(27) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(4)(28) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(4)(29) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(4)(30) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(4)(31) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(4)(32) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(4)(33) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(4)(34) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(4)(35) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(4)(36) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(4)(37) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(4)(38) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(4)(39) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(4)(40) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(4)(41) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(4)(42) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(4)(43) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(4)(44) <= SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1);
SL0_map(4)(45) <= SL0_TSHit(66)(3) or SL0_TSHit(66)(2) or SL0_TSHit(67)(1);
SL0_map(5)(0) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(5)(1) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(5)(2) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(5)(3) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(5)(4) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(5)(5) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(5)(6) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(5)(7) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(5)(8) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(5)(9) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(5)(10) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(5)(11) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(5)(12) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(5)(13) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(5)(14) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(5)(15) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(5)(16) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(5)(17) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(5)(18) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(5)(19) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(5)(20) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(5)(21) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(5)(22) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(5)(23) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(5)(24) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(5)(25) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(5)(26) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(5)(27) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(5)(28) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(5)(29) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(5)(30) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(5)(31) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(5)(32) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(5)(33) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(5)(34) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(5)(35) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(5)(36) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(5)(37) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(5)(38) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(5)(39) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(5)(40) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(5)(41) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(5)(42) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(5)(43) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(5)(44) <= SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1);
SL0_map(5)(45) <= SL0_TSHit(66)(3) or SL0_TSHit(66)(2) or SL0_TSHit(67)(1);
SL0_map(6)(0) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(6)(1) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(6)(2) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(6)(3) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(6)(4) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(6)(5) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(6)(6) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(6)(7) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(6)(8) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(6)(9) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(6)(10) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(6)(11) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(6)(12) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(6)(13) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(6)(14) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(6)(15) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(6)(16) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(6)(17) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(6)(18) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(6)(19) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(6)(20) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(6)(21) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(6)(22) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(6)(23) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(6)(24) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(6)(25) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(6)(26) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(6)(27) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(6)(28) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(6)(29) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(6)(30) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(6)(31) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(6)(32) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(6)(33) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(6)(34) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(6)(35) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(6)(36) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(6)(37) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(6)(38) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(6)(39) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(6)(40) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(6)(41) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(6)(42) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(6)(43) <= SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(6)(44) <= SL0_TSHit(64)(2) or SL0_TSHit(65)(1) or SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1);
SL0_map(6)(45) <= SL0_TSHit(65)(2) or SL0_TSHit(66)(1) or SL0_TSHit(66)(3) or SL0_TSHit(66)(2) or SL0_TSHit(67)(1);
SL0_map(7)(0) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(7)(1) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(7)(2) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(7)(3) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(7)(4) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(7)(5) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(7)(6) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(7)(7) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(7)(8) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(7)(9) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(7)(10) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(7)(11) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(7)(12) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(7)(13) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(7)(14) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(7)(15) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(7)(16) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(7)(17) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(7)(18) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(7)(19) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(7)(20) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(7)(21) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(7)(22) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(7)(23) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(7)(24) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(7)(25) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(7)(26) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(7)(27) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(7)(28) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(7)(29) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(7)(30) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(7)(31) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(7)(32) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(7)(33) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(7)(34) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(7)(35) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(7)(36) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(7)(37) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(7)(38) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(7)(39) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(7)(40) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(7)(41) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(7)(42) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(7)(43) <= SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3);
SL0_map(7)(44) <= SL0_TSHit(64)(2) or SL0_TSHit(65)(1) or SL0_TSHit(65)(3);
SL0_map(7)(45) <= SL0_TSHit(65)(2) or SL0_TSHit(66)(1) or SL0_TSHit(66)(3);
SL0_map(8)(0) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(8)(1) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(8)(2) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(8)(3) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(8)(4) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(8)(5) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(8)(6) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(8)(7) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(8)(8) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(8)(9) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(8)(10) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(8)(11) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(8)(12) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(8)(13) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(8)(14) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(8)(15) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(8)(16) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(8)(17) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(8)(18) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(8)(19) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(8)(20) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(8)(21) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(8)(22) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(8)(23) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(8)(24) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(8)(25) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(8)(26) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(8)(27) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(8)(28) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(8)(29) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(8)(30) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(8)(31) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(8)(32) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(8)(33) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(8)(34) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(8)(35) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(8)(36) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(8)(37) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(8)(38) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(8)(39) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(8)(40) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(8)(41) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(8)(42) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(8)(43) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3);
SL0_map(8)(44) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1) or SL0_TSHit(65)(3);
SL0_map(8)(45) <= SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1) or SL0_TSHit(66)(3);
SL0_map(9)(0) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(9)(1) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(9)(2) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(9)(3) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(9)(4) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(9)(5) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(9)(6) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(9)(7) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(9)(8) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(9)(9) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(9)(10) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(9)(11) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(9)(12) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(9)(13) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(9)(14) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(9)(15) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(9)(16) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(9)(17) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(9)(18) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(9)(19) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(9)(20) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(9)(21) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(9)(22) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(9)(23) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(9)(24) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(9)(25) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(9)(26) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(9)(27) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(9)(28) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(9)(29) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(9)(30) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(9)(31) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(9)(32) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(9)(33) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(9)(34) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(9)(35) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(9)(36) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(9)(37) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(9)(38) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(9)(39) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(9)(40) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(9)(41) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(9)(42) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(9)(43) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(9)(44) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(9)(45) <= SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1);
SL0_map(10)(0) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(10)(1) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(10)(2) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(10)(3) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(10)(4) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(10)(5) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(10)(6) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(10)(7) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(10)(8) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(10)(9) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(10)(10) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(10)(11) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(10)(12) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(10)(13) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(10)(14) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(10)(15) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(10)(16) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(10)(17) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(10)(18) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(10)(19) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(10)(20) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(10)(21) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(10)(22) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(10)(23) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(10)(24) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(10)(25) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(10)(26) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(10)(27) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(10)(28) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(10)(29) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(10)(30) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(10)(31) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(10)(32) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(10)(33) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(10)(34) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(10)(35) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(10)(36) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(10)(37) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(10)(38) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(10)(39) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(10)(40) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(10)(41) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(10)(42) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(10)(43) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(10)(44) <= SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(10)(45) <= SL0_TSHit(64)(2) or SL0_TSHit(65)(1) or SL0_TSHit(65)(3) or SL0_TSHit(65)(2) or SL0_TSHit(66)(1);
SL0_map(11)(0) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(11)(1) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(11)(2) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(11)(3) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(11)(4) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(11)(5) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(11)(6) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(11)(7) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(11)(8) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(11)(9) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(11)(10) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(11)(11) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(11)(12) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(11)(13) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(11)(14) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(11)(15) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(11)(16) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(11)(17) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(11)(18) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(11)(19) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(11)(20) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(11)(21) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(11)(22) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(11)(23) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(11)(24) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(11)(25) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(11)(26) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(11)(27) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(11)(28) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(11)(29) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(11)(30) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(11)(31) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(11)(32) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(11)(33) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(11)(34) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(11)(35) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(11)(36) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(11)(37) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(11)(38) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(11)(39) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(11)(40) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(11)(41) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(11)(42) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(11)(43) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(11)(44) <= SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3);
SL0_map(11)(45) <= SL0_TSHit(64)(2) or SL0_TSHit(65)(1) or SL0_TSHit(65)(3);
SL0_map(12)(0) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(12)(1) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(12)(2) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(12)(3) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(12)(4) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(12)(5) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(12)(6) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(12)(7) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(12)(8) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(12)(9) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(12)(10) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(12)(11) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(12)(12) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(12)(13) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(12)(14) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(12)(15) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(12)(16) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(12)(17) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(12)(18) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(12)(19) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(12)(20) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(12)(21) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(12)(22) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(12)(23) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(12)(24) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(12)(25) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(12)(26) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(12)(27) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(12)(28) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(12)(29) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(12)(30) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(12)(31) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(12)(32) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(12)(33) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(12)(34) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(12)(35) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(12)(36) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(12)(37) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(12)(38) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(12)(39) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(12)(40) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(12)(41) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(12)(42) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(12)(43) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(12)(44) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3);
SL0_map(12)(45) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1) or SL0_TSHit(65)(3);
SL0_map(13)(0) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(13)(1) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(13)(2) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(13)(3) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(13)(4) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(13)(5) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(13)(6) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(13)(7) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(13)(8) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(13)(9) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(13)(10) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(13)(11) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(13)(12) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(13)(13) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(13)(14) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(13)(15) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(13)(16) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(13)(17) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(13)(18) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(13)(19) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(13)(20) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(13)(21) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(13)(22) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(13)(23) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(13)(24) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(13)(25) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(13)(26) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(13)(27) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(13)(28) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(13)(29) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(13)(30) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(13)(31) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(13)(32) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(13)(33) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(13)(34) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(13)(35) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(13)(36) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(13)(37) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(13)(38) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(13)(39) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(13)(40) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(13)(41) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(13)(42) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(13)(43) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(13)(44) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(13)(45) <= SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(14)(0) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(14)(1) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(14)(2) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(14)(3) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(14)(4) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(14)(5) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(14)(6) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(14)(7) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(14)(8) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(14)(9) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(14)(10) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(14)(11) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(14)(12) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(14)(13) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(14)(14) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(14)(15) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(14)(16) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(14)(17) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(14)(18) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(14)(19) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(14)(20) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(14)(21) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(14)(22) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(14)(23) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(14)(24) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(14)(25) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(14)(26) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(14)(27) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(14)(28) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(14)(29) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(14)(30) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(14)(31) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(14)(32) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(14)(33) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(14)(34) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(14)(35) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(14)(36) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(14)(37) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(14)(38) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(14)(39) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(14)(40) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(14)(41) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(14)(42) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(14)(43) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(14)(44) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(14)(45) <= SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3) or SL0_TSHit(64)(2) or SL0_TSHit(65)(1);
SL0_map(15)(0) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(15)(1) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(15)(2) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(15)(3) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(15)(4) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(15)(5) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(15)(6) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(15)(7) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(15)(8) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(15)(9) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(15)(10) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(15)(11) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(15)(12) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(15)(13) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(15)(14) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(15)(15) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(15)(16) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(15)(17) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(15)(18) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(15)(19) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(15)(20) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(15)(21) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(15)(22) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(15)(23) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(15)(24) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(15)(25) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(15)(26) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(15)(27) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(15)(28) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(15)(29) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(15)(30) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(15)(31) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(15)(32) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(15)(33) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(15)(34) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(15)(35) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(15)(36) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(15)(37) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(15)(38) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(15)(39) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(15)(40) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(15)(41) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(15)(42) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(15)(43) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(15)(44) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(15)(45) <= SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3);
SL0_map(16)(0) <= SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(16)(1) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(16)(2) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(16)(3) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(16)(4) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(16)(5) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(16)(6) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(16)(7) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(16)(8) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(16)(9) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(16)(10) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(16)(11) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(16)(12) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(16)(13) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(16)(14) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(16)(15) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(16)(16) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(16)(17) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(16)(18) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(16)(19) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(16)(20) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(16)(21) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(16)(22) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(16)(23) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(16)(24) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(16)(25) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(16)(26) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(16)(27) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(16)(28) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(16)(29) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(16)(30) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(16)(31) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(16)(32) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(16)(33) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(16)(34) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(16)(35) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(16)(36) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(16)(37) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(16)(38) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(16)(39) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(16)(40) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(16)(41) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(16)(42) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(16)(43) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(16)(44) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(16)(45) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3);
SL0_map(17)(0) <= SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(17)(1) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(17)(2) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(17)(3) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(17)(4) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(17)(5) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(17)(6) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(17)(7) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(17)(8) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(17)(9) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(17)(10) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(17)(11) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(17)(12) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(17)(13) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(17)(14) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(17)(15) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(17)(16) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(17)(17) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(17)(18) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(17)(19) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(17)(20) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(17)(21) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(17)(22) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(17)(23) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(17)(24) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(17)(25) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(17)(26) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(17)(27) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(17)(28) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(17)(29) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(17)(30) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(17)(31) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(17)(32) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(17)(33) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(17)(34) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(17)(35) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(17)(36) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(17)(37) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(17)(38) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(17)(39) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(17)(40) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(17)(41) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(17)(42) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(17)(43) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(17)(44) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(17)(45) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1) or SL0_TSHit(64)(3);
SL0_map(18)(0) <= SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1);
SL0_map(18)(1) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(18)(2) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(18)(3) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(18)(4) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(18)(5) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(18)(6) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(18)(7) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(18)(8) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(18)(9) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(18)(10) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(18)(11) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(18)(12) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(18)(13) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(18)(14) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(18)(15) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(18)(16) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(18)(17) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(18)(18) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(18)(19) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(18)(20) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(18)(21) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(18)(22) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(18)(23) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(18)(24) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(18)(25) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(18)(26) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(18)(27) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(18)(28) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(18)(29) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(18)(30) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(18)(31) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(18)(32) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(18)(33) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(18)(34) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(18)(35) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(18)(36) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(18)(37) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(18)(38) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(18)(39) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(18)(40) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(18)(41) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(18)(42) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(18)(43) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(18)(44) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(18)(45) <= SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(19)(0) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1);
SL0_map(19)(1) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(19)(2) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(19)(3) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(19)(4) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(19)(5) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(19)(6) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(19)(7) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(19)(8) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(19)(9) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(19)(10) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(19)(11) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(19)(12) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(19)(13) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(19)(14) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(19)(15) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(19)(16) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(19)(17) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(19)(18) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(19)(19) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(19)(20) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(19)(21) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(19)(22) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(19)(23) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(19)(24) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(19)(25) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(19)(26) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(19)(27) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(19)(28) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(19)(29) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(19)(30) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(19)(31) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(19)(32) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(19)(33) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(19)(34) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(19)(35) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(19)(36) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(19)(37) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(19)(38) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(19)(39) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(19)(40) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(19)(41) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(19)(42) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(19)(43) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(19)(44) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(19)(45) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3) or SL0_TSHit(63)(2) or SL0_TSHit(64)(1);
SL0_map(20)(0) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(20)(1) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(20)(2) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(20)(3) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(20)(4) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(20)(5) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(20)(6) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(20)(7) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(20)(8) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(20)(9) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(20)(10) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(20)(11) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(20)(12) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(20)(13) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(20)(14) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(20)(15) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(20)(16) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(20)(17) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(20)(18) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(20)(19) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(20)(20) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(20)(21) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(20)(22) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(20)(23) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(20)(24) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(20)(25) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(20)(26) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(20)(27) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(20)(28) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(20)(29) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(20)(30) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(20)(31) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(20)(32) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(20)(33) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(20)(34) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(20)(35) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(20)(36) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(20)(37) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(20)(38) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(20)(39) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(20)(40) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(20)(41) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(20)(42) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(20)(43) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(20)(44) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(20)(45) <= SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(21)(0) <= SL0_TSHit(17)(3) or SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(21)(1) <= SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(21)(2) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(21)(3) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(21)(4) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(21)(5) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(21)(6) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(21)(7) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(21)(8) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(21)(9) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(21)(10) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(21)(11) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(21)(12) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(21)(13) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(21)(14) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(21)(15) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(21)(16) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(21)(17) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(21)(18) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(21)(19) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(21)(20) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(21)(21) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(21)(22) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(21)(23) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(21)(24) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(21)(25) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(21)(26) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(21)(27) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(21)(28) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(21)(29) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(21)(30) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(21)(31) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(21)(32) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(21)(33) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(21)(34) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(21)(35) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(21)(36) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(21)(37) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(21)(38) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(21)(39) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(21)(40) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(21)(41) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(21)(42) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(21)(43) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(21)(44) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(21)(45) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1) or SL0_TSHit(63)(3);
SL0_map(22)(0) <= SL0_TSHit(17)(3) or SL0_TSHit(17)(2) or SL0_TSHit(18)(1);
SL0_map(22)(1) <= SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1);
SL0_map(22)(2) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(22)(3) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(22)(4) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(22)(5) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(22)(6) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(22)(7) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(22)(8) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(22)(9) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(22)(10) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(22)(11) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(22)(12) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(22)(13) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(22)(14) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(22)(15) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(22)(16) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(22)(17) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(22)(18) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(22)(19) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(22)(20) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(22)(21) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(22)(22) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(22)(23) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(22)(24) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(22)(25) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(22)(26) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(22)(27) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(22)(28) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(22)(29) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(22)(30) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(22)(31) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(22)(32) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(22)(33) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(22)(34) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(22)(35) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(22)(36) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(22)(37) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(22)(38) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(22)(39) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(22)(40) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(22)(41) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(22)(42) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(22)(43) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(22)(44) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(22)(45) <= SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(23)(0) <= SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3) or SL0_TSHit(17)(2) or SL0_TSHit(18)(1);
SL0_map(23)(1) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1);
SL0_map(23)(2) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(23)(3) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(23)(4) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(23)(5) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(23)(6) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(23)(7) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(23)(8) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(23)(9) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(23)(10) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(23)(11) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(23)(12) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(23)(13) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(23)(14) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(23)(15) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(23)(16) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(23)(17) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(23)(18) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(23)(19) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(23)(20) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(23)(21) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(23)(22) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(23)(23) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(23)(24) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(23)(25) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(23)(26) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(23)(27) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(23)(28) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(23)(29) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(23)(30) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(23)(31) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(23)(32) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(23)(33) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(23)(34) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(23)(35) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(23)(36) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(23)(37) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(23)(38) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(23)(39) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(23)(40) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(23)(41) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(23)(42) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(23)(43) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(23)(44) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(23)(45) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3) or SL0_TSHit(62)(2) or SL0_TSHit(63)(1);
SL0_map(24)(0) <= SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3);
SL0_map(24)(1) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(24)(2) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(24)(3) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(24)(4) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(24)(5) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(24)(6) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(24)(7) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(24)(8) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(24)(9) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(24)(10) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(24)(11) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(24)(12) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(24)(13) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(24)(14) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(24)(15) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(24)(16) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(24)(17) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(24)(18) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(24)(19) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(24)(20) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(24)(21) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(24)(22) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(24)(23) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(24)(24) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(24)(25) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(24)(26) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(24)(27) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(24)(28) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(24)(29) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(24)(30) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(24)(31) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(24)(32) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(24)(33) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(24)(34) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(24)(35) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(24)(36) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(24)(37) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(24)(38) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(24)(39) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(24)(40) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(24)(41) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(24)(42) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(24)(43) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(24)(44) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(24)(45) <= SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(25)(0) <= SL0_TSHit(16)(3) or SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3);
SL0_map(25)(1) <= SL0_TSHit(17)(3) or SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(25)(2) <= SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(25)(3) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(25)(4) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(25)(5) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(25)(6) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(25)(7) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(25)(8) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(25)(9) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(25)(10) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(25)(11) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(25)(12) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(25)(13) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(25)(14) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(25)(15) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(25)(16) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(25)(17) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(25)(18) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(25)(19) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(25)(20) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(25)(21) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(25)(22) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(25)(23) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(25)(24) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(25)(25) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(25)(26) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(25)(27) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(25)(28) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(25)(29) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(25)(30) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(25)(31) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(25)(32) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(25)(33) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(25)(34) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(25)(35) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(25)(36) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(25)(37) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(25)(38) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(25)(39) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(25)(40) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(25)(41) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(25)(42) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(25)(43) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(25)(44) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(25)(45) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1) or SL0_TSHit(62)(3);
SL0_map(26)(0) <= SL0_TSHit(16)(3) or SL0_TSHit(16)(2) or SL0_TSHit(17)(1);
SL0_map(26)(1) <= SL0_TSHit(17)(3) or SL0_TSHit(17)(2) or SL0_TSHit(18)(1);
SL0_map(26)(2) <= SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1);
SL0_map(26)(3) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(26)(4) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(26)(5) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(26)(6) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(26)(7) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(26)(8) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(26)(9) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(26)(10) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(26)(11) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(26)(12) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(26)(13) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(26)(14) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(26)(15) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(26)(16) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(26)(17) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(26)(18) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(26)(19) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(26)(20) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(26)(21) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(26)(22) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(26)(23) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(26)(24) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(26)(25) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(26)(26) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(26)(27) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(26)(28) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(26)(29) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(26)(30) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(26)(31) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(26)(32) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(26)(33) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(26)(34) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(26)(35) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(26)(36) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(26)(37) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(26)(38) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(26)(39) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(26)(40) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(26)(41) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(26)(42) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(26)(43) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(26)(44) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(26)(45) <= SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(27)(0) <= SL0_TSHit(15)(2) or SL0_TSHit(16)(1) or SL0_TSHit(16)(3) or SL0_TSHit(16)(2) or SL0_TSHit(17)(1);
SL0_map(27)(1) <= SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3) or SL0_TSHit(17)(2) or SL0_TSHit(18)(1);
SL0_map(27)(2) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1);
SL0_map(27)(3) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(27)(4) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(27)(5) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(27)(6) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(27)(7) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(27)(8) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(27)(9) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(27)(10) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(27)(11) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(27)(12) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(27)(13) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(27)(14) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(27)(15) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(27)(16) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(27)(17) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(27)(18) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(27)(19) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(27)(20) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(27)(21) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(27)(22) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(27)(23) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(27)(24) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(27)(25) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(27)(26) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(27)(27) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(27)(28) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(27)(29) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(27)(30) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(27)(31) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(27)(32) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(27)(33) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(27)(34) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(27)(35) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(27)(36) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(27)(37) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(27)(38) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(27)(39) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(27)(40) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(27)(41) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(27)(42) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(27)(43) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(27)(44) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(27)(45) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3) or SL0_TSHit(61)(2) or SL0_TSHit(62)(1);
SL0_map(28)(0) <= SL0_TSHit(15)(2) or SL0_TSHit(16)(1) or SL0_TSHit(16)(3);
SL0_map(28)(1) <= SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3);
SL0_map(28)(2) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(28)(3) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(28)(4) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(28)(5) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(28)(6) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(28)(7) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(28)(8) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(28)(9) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(28)(10) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(28)(11) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(28)(12) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(28)(13) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(28)(14) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(28)(15) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(28)(16) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(28)(17) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(28)(18) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(28)(19) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(28)(20) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(28)(21) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(28)(22) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(28)(23) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(28)(24) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(28)(25) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(28)(26) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(28)(27) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(28)(28) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(28)(29) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(28)(30) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(28)(31) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(28)(32) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(28)(33) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(28)(34) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(28)(35) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(28)(36) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(28)(37) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(28)(38) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(28)(39) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(28)(40) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(28)(41) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(28)(42) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(28)(43) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(28)(44) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(28)(45) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(29)(0) <= SL0_TSHit(15)(2) or SL0_TSHit(16)(1) or SL0_TSHit(16)(3);
SL0_map(29)(1) <= SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3);
SL0_map(29)(2) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(29)(3) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(29)(4) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(29)(5) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(29)(6) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(29)(7) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(29)(8) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(29)(9) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(29)(10) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(29)(11) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(29)(12) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(29)(13) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(29)(14) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(29)(15) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(29)(16) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(29)(17) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(29)(18) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(29)(19) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(29)(20) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(29)(21) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(29)(22) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(29)(23) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(29)(24) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(29)(25) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(29)(26) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(29)(27) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(29)(28) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(29)(29) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(29)(30) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(29)(31) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(29)(32) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(29)(33) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(29)(34) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(29)(35) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(29)(36) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(29)(37) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(29)(38) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(29)(39) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(29)(40) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(29)(41) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(29)(42) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(29)(43) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(29)(44) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(29)(45) <= SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(30)(0) <= SL0_TSHit(15)(3) or SL0_TSHit(15)(2) or SL0_TSHit(16)(1) or SL0_TSHit(16)(3);
SL0_map(30)(1) <= SL0_TSHit(16)(3) or SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3);
SL0_map(30)(2) <= SL0_TSHit(17)(3) or SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(30)(3) <= SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(30)(4) <= SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(30)(5) <= SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(30)(6) <= SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(30)(7) <= SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(30)(8) <= SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(30)(9) <= SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(30)(10) <= SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(30)(11) <= SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(30)(12) <= SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(30)(13) <= SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(30)(14) <= SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(30)(15) <= SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(30)(16) <= SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(30)(17) <= SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(30)(18) <= SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(30)(19) <= SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(30)(20) <= SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(30)(21) <= SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(30)(22) <= SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(30)(23) <= SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(30)(24) <= SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(30)(25) <= SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(30)(26) <= SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(30)(27) <= SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(30)(28) <= SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(30)(29) <= SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(30)(30) <= SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(30)(31) <= SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(30)(32) <= SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(30)(33) <= SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(30)(34) <= SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(30)(35) <= SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(30)(36) <= SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(30)(37) <= SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(30)(38) <= SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(30)(39) <= SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(30)(40) <= SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(30)(41) <= SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(30)(42) <= SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(30)(43) <= SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(30)(44) <= SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(30)(45) <= SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1) or SL0_TSHit(61)(3);
SL0_map(31)(0) <= SL0_TSHit(14)(2) or SL0_TSHit(15)(1) or SL0_TSHit(15)(3) or SL0_TSHit(15)(2) or SL0_TSHit(16)(1);
SL0_map(31)(1) <= SL0_TSHit(15)(2) or SL0_TSHit(16)(1) or SL0_TSHit(16)(3) or SL0_TSHit(16)(2) or SL0_TSHit(17)(1);
SL0_map(31)(2) <= SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3) or SL0_TSHit(17)(2) or SL0_TSHit(18)(1);
SL0_map(31)(3) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3) or SL0_TSHit(18)(2) or SL0_TSHit(19)(1);
SL0_map(31)(4) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3) or SL0_TSHit(19)(2) or SL0_TSHit(20)(1);
SL0_map(31)(5) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3) or SL0_TSHit(20)(2) or SL0_TSHit(21)(1);
SL0_map(31)(6) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3) or SL0_TSHit(21)(2) or SL0_TSHit(22)(1);
SL0_map(31)(7) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3) or SL0_TSHit(22)(2) or SL0_TSHit(23)(1);
SL0_map(31)(8) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3) or SL0_TSHit(23)(2) or SL0_TSHit(24)(1);
SL0_map(31)(9) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3) or SL0_TSHit(24)(2) or SL0_TSHit(25)(1);
SL0_map(31)(10) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3) or SL0_TSHit(25)(2) or SL0_TSHit(26)(1);
SL0_map(31)(11) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3) or SL0_TSHit(26)(2) or SL0_TSHit(27)(1);
SL0_map(31)(12) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3) or SL0_TSHit(27)(2) or SL0_TSHit(28)(1);
SL0_map(31)(13) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3) or SL0_TSHit(28)(2) or SL0_TSHit(29)(1);
SL0_map(31)(14) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3) or SL0_TSHit(29)(2) or SL0_TSHit(30)(1);
SL0_map(31)(15) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3) or SL0_TSHit(30)(2) or SL0_TSHit(31)(1);
SL0_map(31)(16) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3) or SL0_TSHit(31)(2) or SL0_TSHit(32)(1);
SL0_map(31)(17) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3) or SL0_TSHit(32)(2) or SL0_TSHit(33)(1);
SL0_map(31)(18) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3) or SL0_TSHit(33)(2) or SL0_TSHit(34)(1);
SL0_map(31)(19) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3) or SL0_TSHit(34)(2) or SL0_TSHit(35)(1);
SL0_map(31)(20) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3) or SL0_TSHit(35)(2) or SL0_TSHit(36)(1);
SL0_map(31)(21) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3) or SL0_TSHit(36)(2) or SL0_TSHit(37)(1);
SL0_map(31)(22) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3) or SL0_TSHit(37)(2) or SL0_TSHit(38)(1);
SL0_map(31)(23) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3) or SL0_TSHit(38)(2) or SL0_TSHit(39)(1);
SL0_map(31)(24) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3) or SL0_TSHit(39)(2) or SL0_TSHit(40)(1);
SL0_map(31)(25) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3) or SL0_TSHit(40)(2) or SL0_TSHit(41)(1);
SL0_map(31)(26) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3) or SL0_TSHit(41)(2) or SL0_TSHit(42)(1);
SL0_map(31)(27) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3) or SL0_TSHit(42)(2) or SL0_TSHit(43)(1);
SL0_map(31)(28) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3) or SL0_TSHit(43)(2) or SL0_TSHit(44)(1);
SL0_map(31)(29) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3) or SL0_TSHit(44)(2) or SL0_TSHit(45)(1);
SL0_map(31)(30) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3) or SL0_TSHit(45)(2) or SL0_TSHit(46)(1);
SL0_map(31)(31) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3) or SL0_TSHit(46)(2) or SL0_TSHit(47)(1);
SL0_map(31)(32) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3) or SL0_TSHit(47)(2) or SL0_TSHit(48)(1);
SL0_map(31)(33) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3) or SL0_TSHit(48)(2) or SL0_TSHit(49)(1);
SL0_map(31)(34) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3) or SL0_TSHit(49)(2) or SL0_TSHit(50)(1);
SL0_map(31)(35) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3) or SL0_TSHit(50)(2) or SL0_TSHit(51)(1);
SL0_map(31)(36) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3) or SL0_TSHit(51)(2) or SL0_TSHit(52)(1);
SL0_map(31)(37) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3) or SL0_TSHit(52)(2) or SL0_TSHit(53)(1);
SL0_map(31)(38) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3) or SL0_TSHit(53)(2) or SL0_TSHit(54)(1);
SL0_map(31)(39) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3) or SL0_TSHit(54)(2) or SL0_TSHit(55)(1);
SL0_map(31)(40) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3) or SL0_TSHit(55)(2) or SL0_TSHit(56)(1);
SL0_map(31)(41) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3) or SL0_TSHit(56)(2) or SL0_TSHit(57)(1);
SL0_map(31)(42) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3) or SL0_TSHit(57)(2) or SL0_TSHit(58)(1);
SL0_map(31)(43) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3) or SL0_TSHit(58)(2) or SL0_TSHit(59)(1);
SL0_map(31)(44) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3) or SL0_TSHit(59)(2) or SL0_TSHit(60)(1);
SL0_map(31)(45) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3) or SL0_TSHit(60)(2) or SL0_TSHit(61)(1);
SL0_map(32)(0) <= SL0_TSHit(14)(2) or SL0_TSHit(15)(1) or SL0_TSHit(15)(3);
SL0_map(32)(1) <= SL0_TSHit(15)(2) or SL0_TSHit(16)(1) or SL0_TSHit(16)(3);
SL0_map(32)(2) <= SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3);
SL0_map(32)(3) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(32)(4) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(32)(5) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(32)(6) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(32)(7) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(32)(8) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(32)(9) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(32)(10) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(32)(11) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(32)(12) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(32)(13) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(32)(14) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(32)(15) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(32)(16) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(32)(17) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(32)(18) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(32)(19) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(32)(20) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(32)(21) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(32)(22) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(32)(23) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(32)(24) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(32)(25) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(32)(26) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(32)(27) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(32)(28) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(32)(29) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(32)(30) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(32)(31) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(32)(32) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(32)(33) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(32)(34) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(32)(35) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(32)(36) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(32)(37) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(32)(38) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(32)(39) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(32)(40) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(32)(41) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(32)(42) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(32)(43) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(32)(44) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(32)(45) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
SL0_map(33)(0) <= SL0_TSHit(14)(2) or SL0_TSHit(15)(1) or SL0_TSHit(15)(3);
SL0_map(33)(1) <= SL0_TSHit(15)(2) or SL0_TSHit(16)(1) or SL0_TSHit(16)(3);
SL0_map(33)(2) <= SL0_TSHit(16)(2) or SL0_TSHit(17)(1) or SL0_TSHit(17)(3);
SL0_map(33)(3) <= SL0_TSHit(17)(2) or SL0_TSHit(18)(1) or SL0_TSHit(18)(3);
SL0_map(33)(4) <= SL0_TSHit(18)(2) or SL0_TSHit(19)(1) or SL0_TSHit(19)(3);
SL0_map(33)(5) <= SL0_TSHit(19)(2) or SL0_TSHit(20)(1) or SL0_TSHit(20)(3);
SL0_map(33)(6) <= SL0_TSHit(20)(2) or SL0_TSHit(21)(1) or SL0_TSHit(21)(3);
SL0_map(33)(7) <= SL0_TSHit(21)(2) or SL0_TSHit(22)(1) or SL0_TSHit(22)(3);
SL0_map(33)(8) <= SL0_TSHit(22)(2) or SL0_TSHit(23)(1) or SL0_TSHit(23)(3);
SL0_map(33)(9) <= SL0_TSHit(23)(2) or SL0_TSHit(24)(1) or SL0_TSHit(24)(3);
SL0_map(33)(10) <= SL0_TSHit(24)(2) or SL0_TSHit(25)(1) or SL0_TSHit(25)(3);
SL0_map(33)(11) <= SL0_TSHit(25)(2) or SL0_TSHit(26)(1) or SL0_TSHit(26)(3);
SL0_map(33)(12) <= SL0_TSHit(26)(2) or SL0_TSHit(27)(1) or SL0_TSHit(27)(3);
SL0_map(33)(13) <= SL0_TSHit(27)(2) or SL0_TSHit(28)(1) or SL0_TSHit(28)(3);
SL0_map(33)(14) <= SL0_TSHit(28)(2) or SL0_TSHit(29)(1) or SL0_TSHit(29)(3);
SL0_map(33)(15) <= SL0_TSHit(29)(2) or SL0_TSHit(30)(1) or SL0_TSHit(30)(3);
SL0_map(33)(16) <= SL0_TSHit(30)(2) or SL0_TSHit(31)(1) or SL0_TSHit(31)(3);
SL0_map(33)(17) <= SL0_TSHit(31)(2) or SL0_TSHit(32)(1) or SL0_TSHit(32)(3);
SL0_map(33)(18) <= SL0_TSHit(32)(2) or SL0_TSHit(33)(1) or SL0_TSHit(33)(3);
SL0_map(33)(19) <= SL0_TSHit(33)(2) or SL0_TSHit(34)(1) or SL0_TSHit(34)(3);
SL0_map(33)(20) <= SL0_TSHit(34)(2) or SL0_TSHit(35)(1) or SL0_TSHit(35)(3);
SL0_map(33)(21) <= SL0_TSHit(35)(2) or SL0_TSHit(36)(1) or SL0_TSHit(36)(3);
SL0_map(33)(22) <= SL0_TSHit(36)(2) or SL0_TSHit(37)(1) or SL0_TSHit(37)(3);
SL0_map(33)(23) <= SL0_TSHit(37)(2) or SL0_TSHit(38)(1) or SL0_TSHit(38)(3);
SL0_map(33)(24) <= SL0_TSHit(38)(2) or SL0_TSHit(39)(1) or SL0_TSHit(39)(3);
SL0_map(33)(25) <= SL0_TSHit(39)(2) or SL0_TSHit(40)(1) or SL0_TSHit(40)(3);
SL0_map(33)(26) <= SL0_TSHit(40)(2) or SL0_TSHit(41)(1) or SL0_TSHit(41)(3);
SL0_map(33)(27) <= SL0_TSHit(41)(2) or SL0_TSHit(42)(1) or SL0_TSHit(42)(3);
SL0_map(33)(28) <= SL0_TSHit(42)(2) or SL0_TSHit(43)(1) or SL0_TSHit(43)(3);
SL0_map(33)(29) <= SL0_TSHit(43)(2) or SL0_TSHit(44)(1) or SL0_TSHit(44)(3);
SL0_map(33)(30) <= SL0_TSHit(44)(2) or SL0_TSHit(45)(1) or SL0_TSHit(45)(3);
SL0_map(33)(31) <= SL0_TSHit(45)(2) or SL0_TSHit(46)(1) or SL0_TSHit(46)(3);
SL0_map(33)(32) <= SL0_TSHit(46)(2) or SL0_TSHit(47)(1) or SL0_TSHit(47)(3);
SL0_map(33)(33) <= SL0_TSHit(47)(2) or SL0_TSHit(48)(1) or SL0_TSHit(48)(3);
SL0_map(33)(34) <= SL0_TSHit(48)(2) or SL0_TSHit(49)(1) or SL0_TSHit(49)(3);
SL0_map(33)(35) <= SL0_TSHit(49)(2) or SL0_TSHit(50)(1) or SL0_TSHit(50)(3);
SL0_map(33)(36) <= SL0_TSHit(50)(2) or SL0_TSHit(51)(1) or SL0_TSHit(51)(3);
SL0_map(33)(37) <= SL0_TSHit(51)(2) or SL0_TSHit(52)(1) or SL0_TSHit(52)(3);
SL0_map(33)(38) <= SL0_TSHit(52)(2) or SL0_TSHit(53)(1) or SL0_TSHit(53)(3);
SL0_map(33)(39) <= SL0_TSHit(53)(2) or SL0_TSHit(54)(1) or SL0_TSHit(54)(3);
SL0_map(33)(40) <= SL0_TSHit(54)(2) or SL0_TSHit(55)(1) or SL0_TSHit(55)(3);
SL0_map(33)(41) <= SL0_TSHit(55)(2) or SL0_TSHit(56)(1) or SL0_TSHit(56)(3);
SL0_map(33)(42) <= SL0_TSHit(56)(2) or SL0_TSHit(57)(1) or SL0_TSHit(57)(3);
SL0_map(33)(43) <= SL0_TSHit(57)(2) or SL0_TSHit(58)(1) or SL0_TSHit(58)(3);
SL0_map(33)(44) <= SL0_TSHit(58)(2) or SL0_TSHit(59)(1) or SL0_TSHit(59)(3);
SL0_map(33)(45) <= SL0_TSHit(59)(2) or SL0_TSHit(60)(1) or SL0_TSHit(60)(3);
 
end Behavioral;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
 
entity UT3_0_SL8_P is
 
Port (
           SL8_row1  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row2  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row3  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row4  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row5  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row6  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row7  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row8  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row9  : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row10 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row11 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row12 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row13 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row14 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row15 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_row16 : out  STD_LOGIC_VECTOR (39 downto 0);
           SL8_TS    : in   STD_LOGIC_VECTOR (192 downto 0));
end UT3_0_SL8_P;
 
 
architecture Behavioral of UT3_0_SL8_P is
 
begin
 
SL8_row1(0)<=SL8_TS(41) or SL8_TS(42) or SL8_TS(43) or SL8_TS(44) or SL8_TS(45) or SL8_TS(46) or SL8_TS(47) or SL8_TS(48) or SL8_TS(49) or SL8_TS(50) or SL8_TS(51) or SL8_TS(52) or SL8_TS(53) or SL8_TS(54) or SL8_TS(55) ;
SL8_row1(1)<=SL8_TS(43) or SL8_TS(44) or SL8_TS(45) or SL8_TS(46) or SL8_TS(47) or SL8_TS(48) or SL8_TS(49) or SL8_TS(50) or SL8_TS(51) or SL8_TS(52) or SL8_TS(53) or SL8_TS(54) or SL8_TS(55) or SL8_TS(56) or SL8_TS(57) ;
SL8_row1(2)<=SL8_TS(45) or SL8_TS(46) or SL8_TS(47) or SL8_TS(48) or SL8_TS(49) or SL8_TS(50) or SL8_TS(51) or SL8_TS(52) or SL8_TS(53) or SL8_TS(54) or SL8_TS(55) or SL8_TS(56) or SL8_TS(57) or SL8_TS(58) or SL8_TS(59) ;
SL8_row1(3)<=SL8_TS(48) or SL8_TS(49) or SL8_TS(50) or SL8_TS(51) or SL8_TS(52) or SL8_TS(53) or SL8_TS(54) or SL8_TS(55) or SL8_TS(56) or SL8_TS(57) or SL8_TS(58) or SL8_TS(59) or SL8_TS(60) or SL8_TS(61) or SL8_TS(62) ;
SL8_row1(4)<=SL8_TS(50) or SL8_TS(51) or SL8_TS(52) or SL8_TS(53) or SL8_TS(54) or SL8_TS(55) or SL8_TS(56) or SL8_TS(57) or SL8_TS(58) or SL8_TS(59) or SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) ;
SL8_row1(5)<=SL8_TS(53) or SL8_TS(54) or SL8_TS(55) or SL8_TS(56) or SL8_TS(57) or SL8_TS(58) or SL8_TS(59) or SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) ;
SL8_row1(6)<=SL8_TS(55) or SL8_TS(56) or SL8_TS(57) or SL8_TS(58) or SL8_TS(59) or SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) ;
SL8_row1(7)<=SL8_TS(57) or SL8_TS(58) or SL8_TS(59) or SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) ;
SL8_row1(8)<=SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) ;
SL8_row1(9)<=SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) ;
SL8_row1(10)<=SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) ;
SL8_row1(11)<=SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) ;
SL8_row1(12)<=SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) ;
SL8_row1(13)<=SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) ;
SL8_row1(14)<=SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) ;
SL8_row1(15)<=SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) ;
SL8_row1(16)<=SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) ;
SL8_row1(17)<=SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row1(18)<=SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) ;
SL8_row1(19)<=SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row1(20)<=SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) ;
SL8_row1(21)<=SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) ;
SL8_row1(22)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row1(23)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) ;
SL8_row1(24)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row1(25)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) ;
SL8_row1(26)<=SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) ;
SL8_row1(27)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row1(28)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) ;
SL8_row1(29)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row1(30)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) ;
SL8_row1(31)<=SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) ;
SL8_row1(32)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row1(33)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) ;
SL8_row1(34)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row1(35)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) ;
SL8_row1(36)<=SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) ;
SL8_row1(37)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row1(38)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) ;
SL8_row1(39)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row2(0)<=SL8_TS(53) or SL8_TS(54) or SL8_TS(55) or SL8_TS(56) or SL8_TS(57) or SL8_TS(58) or SL8_TS(59) or SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) ;
SL8_row2(1)<=SL8_TS(56) or SL8_TS(57) or SL8_TS(58) or SL8_TS(59) or SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) ;
SL8_row2(2)<=SL8_TS(58) or SL8_TS(59) or SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) ;
SL8_row2(3)<=SL8_TS(60) or SL8_TS(61) or SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) ;
SL8_row2(4)<=SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) ;
SL8_row2(5)<=SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) ;
SL8_row2(6)<=SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) ;
SL8_row2(7)<=SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) ;
SL8_row2(8)<=SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) ;
SL8_row2(9)<=SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) ;
SL8_row2(10)<=SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) ;
SL8_row2(11)<=SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) ;
SL8_row2(12)<=SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) ;
SL8_row2(13)<=SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row2(14)<=SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) ;
SL8_row2(15)<=SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row2(16)<=SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) ;
SL8_row2(17)<=SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) ;
SL8_row2(18)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row2(19)<=SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) ;
SL8_row2(20)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row2(21)<=SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) ;
SL8_row2(22)<=SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) ;
SL8_row2(23)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row2(24)<=SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) ;
SL8_row2(25)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row2(26)<=SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) ;
SL8_row2(27)<=SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) ;
SL8_row2(28)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row2(29)<=SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) ;
SL8_row2(30)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row2(31)<=SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) ;
SL8_row2(32)<=SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) ;
SL8_row2(33)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row2(34)<=SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) ;
SL8_row2(35)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row2(36)<=SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) ;
SL8_row2(37)<=SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) ;
SL8_row2(38)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row2(39)<=SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) ;
SL8_row3(0)<=SL8_TS(62) or SL8_TS(63) or SL8_TS(64) or SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) ;
SL8_row3(1)<=SL8_TS(65) or SL8_TS(66) or SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) ;
SL8_row3(2)<=SL8_TS(67) or SL8_TS(68) or SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) ;
SL8_row3(3)<=SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) ;
SL8_row3(4)<=SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) ;
SL8_row3(5)<=SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) ;
SL8_row3(6)<=SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) ;
SL8_row3(7)<=SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) ;
SL8_row3(8)<=SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) ;
SL8_row3(9)<=SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) ;
SL8_row3(10)<=SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) ;
SL8_row3(11)<=SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) ;
SL8_row3(12)<=SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) ;
SL8_row3(13)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) ;
SL8_row3(14)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) ;
SL8_row3(15)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) ;
SL8_row3(16)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) ;
SL8_row3(17)<=SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) ;
SL8_row3(18)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) ;
SL8_row3(19)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) ;
SL8_row3(20)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) ;
SL8_row3(21)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) ;
SL8_row3(22)<=SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) ;
SL8_row3(23)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) ;
SL8_row3(24)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) ;
SL8_row3(25)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) ;
SL8_row3(26)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) ;
SL8_row3(27)<=SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) ;
SL8_row3(28)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) ;
SL8_row3(29)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) ;
SL8_row3(30)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) ;
SL8_row3(31)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) ;
SL8_row3(32)<=SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) ;
SL8_row3(33)<=SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) ;
SL8_row3(34)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) ;
SL8_row3(35)<=SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) ;
SL8_row3(36)<=SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) ;
SL8_row3(37)<=SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) ;
SL8_row3(38)<=SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) ;
SL8_row3(39)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) ;
SL8_row4(0)<=SL8_TS(69) or SL8_TS(70) or SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) ;
SL8_row4(1)<=SL8_TS(71) or SL8_TS(72) or SL8_TS(73) or SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) ;
SL8_row4(2)<=SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) ;
SL8_row4(3)<=SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) ;
SL8_row4(4)<=SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) ;
SL8_row4(5)<=SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) ;
SL8_row4(6)<=SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) ;
SL8_row4(7)<=SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) ;
SL8_row4(8)<=SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row4(9)<=SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) ;
SL8_row4(10)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row4(11)<=SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) ;
SL8_row4(12)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) ;
SL8_row4(13)<=SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row4(14)<=SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) ;
SL8_row4(15)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row4(16)<=SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) ;
SL8_row4(17)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) ;
SL8_row4(18)<=SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row4(19)<=SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) ;
SL8_row4(20)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row4(21)<=SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) ;
SL8_row4(22)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) ;
SL8_row4(23)<=SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row4(24)<=SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) ;
SL8_row4(25)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row4(26)<=SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) ;
SL8_row4(27)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) ;
SL8_row4(28)<=SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row4(29)<=SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) ;
SL8_row4(30)<=SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row4(31)<=SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) ;
SL8_row4(32)<=SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) ;
SL8_row4(33)<=SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row4(34)<=SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) ;
SL8_row4(35)<=SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) ;
SL8_row4(36)<=SL8_TS(155) or SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) ;
SL8_row4(37)<=SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) ;
SL8_row4(38)<=SL8_TS(160) or SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) or SL8_TS(165) or SL8_TS(166) or SL8_TS(167) ;
SL8_row4(39)<=SL8_TS(162) or SL8_TS(163) or SL8_TS(164) or SL8_TS(165) or SL8_TS(166) or SL8_TS(167) or SL8_TS(168) or SL8_TS(169) ;
SL8_row5(0)<=SL8_TS(74) or SL8_TS(75) or SL8_TS(76) or SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) ;
SL8_row5(1)<=SL8_TS(77) or SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) ;
SL8_row5(2)<=SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) ;
SL8_row5(3)<=SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) ;
SL8_row5(4)<=SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) ;
SL8_row5(5)<=SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) ;
SL8_row5(6)<=SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) ;
SL8_row5(7)<=SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) ;
SL8_row5(8)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) ;
SL8_row5(9)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) ;
SL8_row5(10)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) ;
SL8_row5(11)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) ;
SL8_row5(12)<=SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) ;
SL8_row5(13)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) ;
SL8_row5(14)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) ;
SL8_row5(15)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) ;
SL8_row5(16)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) ;
SL8_row5(17)<=SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) ;
SL8_row5(18)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) ;
SL8_row5(19)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) ;
SL8_row5(20)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) ;
SL8_row5(21)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) ;
SL8_row5(22)<=SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) ;
SL8_row5(23)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) ;
SL8_row5(24)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) ;
SL8_row5(25)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) ;
SL8_row5(26)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) ;
SL8_row5(27)<=SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) ;
SL8_row5(28)<=SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) ;
SL8_row5(29)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) ;
SL8_row5(30)<=SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) ;
SL8_row5(31)<=SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) ;
SL8_row5(32)<=SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) ;
SL8_row5(33)<=SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) ;
SL8_row5(34)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) ;
SL8_row5(35)<=SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) ;
SL8_row5(36)<=SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) or SL8_TS(165) or SL8_TS(166) ;
SL8_row5(37)<=SL8_TS(163) or SL8_TS(164) or SL8_TS(165) or SL8_TS(166) or SL8_TS(167) or SL8_TS(168) ;
SL8_row5(38)<=SL8_TS(165) or SL8_TS(166) or SL8_TS(167) or SL8_TS(168) or SL8_TS(169) or SL8_TS(170) or SL8_TS(171) ;
SL8_row5(39)<=SL8_TS(168) or SL8_TS(169) or SL8_TS(170) or SL8_TS(171) or SL8_TS(172) or SL8_TS(173) ;
SL8_row6(0)<=SL8_TS(78) or SL8_TS(79) or SL8_TS(80) or SL8_TS(81) or SL8_TS(82) or SL8_TS(83) ;
SL8_row6(1)<=SL8_TS(81) or SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) ;
SL8_row6(2)<=SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) ;
SL8_row6(3)<=SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) ;
SL8_row6(4)<=SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) ;
SL8_row6(5)<=SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row6(6)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) ;
SL8_row6(7)<=SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row6(8)<=SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) ;
SL8_row6(9)<=SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) ;
SL8_row6(10)<=SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row6(11)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) ;
SL8_row6(12)<=SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row6(13)<=SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) ;
SL8_row6(14)<=SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) ;
SL8_row6(15)<=SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row6(16)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) ;
SL8_row6(17)<=SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row6(18)<=SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) ;
SL8_row6(19)<=SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) ;
SL8_row6(20)<=SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row6(21)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) ;
SL8_row6(22)<=SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row6(23)<=SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) ;
SL8_row6(24)<=SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) ;
SL8_row6(25)<=SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row6(26)<=SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) ;
SL8_row6(27)<=SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row6(28)<=SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) ;
SL8_row6(29)<=SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) ;
SL8_row6(30)<=SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row6(31)<=SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) ;
SL8_row6(32)<=SL8_TS(155) or SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) ;
SL8_row6(33)<=SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) ;
SL8_row6(34)<=SL8_TS(160) or SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) or SL8_TS(165) ;
SL8_row6(35)<=SL8_TS(162) or SL8_TS(163) or SL8_TS(164) or SL8_TS(165) or SL8_TS(166) or SL8_TS(167) ;
SL8_row6(36)<=SL8_TS(165) or SL8_TS(166) or SL8_TS(167) or SL8_TS(168) or SL8_TS(169) ;
SL8_row6(37)<=SL8_TS(167) or SL8_TS(168) or SL8_TS(169) or SL8_TS(170) or SL8_TS(171) or SL8_TS(172) ;
SL8_row6(38)<=SL8_TS(169) or SL8_TS(170) or SL8_TS(171) or SL8_TS(172) or SL8_TS(173) or SL8_TS(174) ;
SL8_row6(39)<=SL8_TS(172) or SL8_TS(173) or SL8_TS(174) or SL8_TS(175) or SL8_TS(176) or SL8_TS(177) ;
SL8_row7(0)<=SL8_TS(82) or SL8_TS(83) or SL8_TS(84) or SL8_TS(85) or SL8_TS(86) ;
SL8_row7(1)<=SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) ;
SL8_row7(2)<=SL8_TS(86) or SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) ;
SL8_row7(3)<=SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) ;
SL8_row7(4)<=SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row7(5)<=SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) ;
SL8_row7(6)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row7(7)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) ;
SL8_row7(8)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) ;
SL8_row7(9)<=SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row7(10)<=SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) ;
SL8_row7(11)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row7(12)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) ;
SL8_row7(13)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) ;
SL8_row7(14)<=SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row7(15)<=SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) ;
SL8_row7(16)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row7(17)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) ;
SL8_row7(18)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) ;
SL8_row7(19)<=SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row7(20)<=SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) ;
SL8_row7(21)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row7(22)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) ;
SL8_row7(23)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) ;
SL8_row7(24)<=SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row7(25)<=SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) ;
SL8_row7(26)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row7(27)<=SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) ;
SL8_row7(28)<=SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) ;
SL8_row7(29)<=SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row7(30)<=SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) or SL8_TS(158) ;
SL8_row7(31)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) ;
SL8_row7(32)<=SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) or SL8_TS(163) ;
SL8_row7(33)<=SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) or SL8_TS(165) ;
SL8_row7(34)<=SL8_TS(163) or SL8_TS(164) or SL8_TS(165) or SL8_TS(166) or SL8_TS(167) ;
SL8_row7(35)<=SL8_TS(166) or SL8_TS(167) or SL8_TS(168) or SL8_TS(169) or SL8_TS(170) ;
SL8_row7(36)<=SL8_TS(168) or SL8_TS(169) or SL8_TS(170) or SL8_TS(171) or SL8_TS(172) ;
SL8_row7(37)<=SL8_TS(170) or SL8_TS(171) or SL8_TS(172) or SL8_TS(173) or SL8_TS(174) or SL8_TS(175) ;
SL8_row7(38)<=SL8_TS(173) or SL8_TS(174) or SL8_TS(175) or SL8_TS(176) or SL8_TS(177) ;
SL8_row7(39)<=SL8_TS(175) or SL8_TS(176) or SL8_TS(177) or SL8_TS(178) or SL8_TS(179) ;
SL8_row8(0)<=SL8_TS(84) or SL8_TS(85) or SL8_TS(86) or SL8_TS(87) or SL8_TS(88) ;
SL8_row8(1)<=SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) ;
SL8_row8(2)<=SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) or SL8_TS(93) ;
SL8_row8(3)<=SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row8(4)<=SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) or SL8_TS(98) ;
SL8_row8(5)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row8(6)<=SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) ;
SL8_row8(7)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) or SL8_TS(105) ;
SL8_row8(8)<=SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row8(9)<=SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) or SL8_TS(110) ;
SL8_row8(10)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row8(11)<=SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) ;
SL8_row8(12)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) or SL8_TS(117) ;
SL8_row8(13)<=SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row8(14)<=SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) or SL8_TS(122) ;
SL8_row8(15)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row8(16)<=SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) ;
SL8_row8(17)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) or SL8_TS(129) ;
SL8_row8(18)<=SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row8(19)<=SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) or SL8_TS(134) ;
SL8_row8(20)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row8(21)<=SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) ;
SL8_row8(22)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) or SL8_TS(141) ;
SL8_row8(23)<=SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row8(24)<=SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) or SL8_TS(146) ;
SL8_row8(25)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row8(26)<=SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) ;
SL8_row8(27)<=SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) or SL8_TS(153) ;
SL8_row8(28)<=SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row8(29)<=SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) or SL8_TS(158) ;
SL8_row8(30)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) ;
SL8_row8(31)<=SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) ;
SL8_row8(32)<=SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) or SL8_TS(165) ;
SL8_row8(33)<=SL8_TS(164) or SL8_TS(165) or SL8_TS(166) or SL8_TS(167) ;
SL8_row8(34)<=SL8_TS(166) or SL8_TS(167) or SL8_TS(168) or SL8_TS(169) or SL8_TS(170) ;
SL8_row8(35)<=SL8_TS(168) or SL8_TS(169) or SL8_TS(170) or SL8_TS(171) or SL8_TS(172) ;
SL8_row8(36)<=SL8_TS(171) or SL8_TS(172) or SL8_TS(173) or SL8_TS(174) ;
SL8_row8(37)<=SL8_TS(173) or SL8_TS(174) or SL8_TS(175) or SL8_TS(176) or SL8_TS(177) ;
SL8_row8(38)<=SL8_TS(176) or SL8_TS(177) or SL8_TS(178) or SL8_TS(179) ;
SL8_row8(39)<=SL8_TS(178) or SL8_TS(179) or SL8_TS(180) or SL8_TS(181) or SL8_TS(182) ;
SL8_row9(0)<=SL8_TS(87) or SL8_TS(88) or SL8_TS(89) or SL8_TS(90) ;
SL8_row9(1)<=SL8_TS(89) or SL8_TS(90) or SL8_TS(91) or SL8_TS(92) ;
SL8_row9(2)<=SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row9(3)<=SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) ;
SL8_row9(4)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) or SL8_TS(99) ;
SL8_row9(5)<=SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) ;
SL8_row9(6)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) or SL8_TS(104) ;
SL8_row9(7)<=SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row9(8)<=SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) ;
SL8_row9(9)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) or SL8_TS(111) ;
SL8_row9(10)<=SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) ;
SL8_row9(11)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) or SL8_TS(116) ;
SL8_row9(12)<=SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row9(13)<=SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) ;
SL8_row9(14)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) or SL8_TS(123) ;
SL8_row9(15)<=SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) ;
SL8_row9(16)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) or SL8_TS(128) ;
SL8_row9(17)<=SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row9(18)<=SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) ;
SL8_row9(19)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) or SL8_TS(135) ;
SL8_row9(20)<=SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) ;
SL8_row9(21)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) or SL8_TS(140) ;
SL8_row9(22)<=SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row9(23)<=SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) ;
SL8_row9(24)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) or SL8_TS(147) ;
SL8_row9(25)<=SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) ;
SL8_row9(26)<=SL8_TS(149) or SL8_TS(150) or SL8_TS(151) or SL8_TS(152) ;
SL8_row9(27)<=SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row9(28)<=SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) ;
SL8_row9(29)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) or SL8_TS(159) ;
SL8_row9(30)<=SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) ;
SL8_row9(31)<=SL8_TS(161) or SL8_TS(162) or SL8_TS(163) or SL8_TS(164) ;
SL8_row9(32)<=SL8_TS(163) or SL8_TS(164) or SL8_TS(165) or SL8_TS(166) or SL8_TS(167) ;
SL8_row9(33)<=SL8_TS(166) or SL8_TS(167) or SL8_TS(168) or SL8_TS(169) ;
SL8_row9(34)<=SL8_TS(168) or SL8_TS(169) or SL8_TS(170) or SL8_TS(171) ;
SL8_row9(35)<=SL8_TS(171) or SL8_TS(172) or SL8_TS(173) or SL8_TS(174) ;
SL8_row9(36)<=SL8_TS(173) or SL8_TS(174) or SL8_TS(175) or SL8_TS(176) ;
SL8_row9(37)<=SL8_TS(175) or SL8_TS(176) or SL8_TS(177) or SL8_TS(178) or SL8_TS(179) ;
SL8_row9(38)<=SL8_TS(178) or SL8_TS(179) or SL8_TS(180) or SL8_TS(181) ;
SL8_row9(39)<=SL8_TS(180) or SL8_TS(181) or SL8_TS(182) or SL8_TS(183) ;
SL8_row10(0)<=SL8_TS(88) or SL8_TS(89) or SL8_TS(90) or SL8_TS(91) ;
SL8_row10(1)<=SL8_TS(91) or SL8_TS(92) or SL8_TS(93) or SL8_TS(94) ;
SL8_row10(2)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) ;
SL8_row10(3)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) ;
SL8_row10(4)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) ;
SL8_row10(5)<=SL8_TS(100) or SL8_TS(101) or SL8_TS(102) or SL8_TS(103) ;
SL8_row10(6)<=SL8_TS(103) or SL8_TS(104) or SL8_TS(105) or SL8_TS(106) ;
SL8_row10(7)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) ;
SL8_row10(8)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) ;
SL8_row10(9)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) ;
SL8_row10(10)<=SL8_TS(112) or SL8_TS(113) or SL8_TS(114) or SL8_TS(115) ;
SL8_row10(11)<=SL8_TS(115) or SL8_TS(116) or SL8_TS(117) or SL8_TS(118) ;
SL8_row10(12)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) ;
SL8_row10(13)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) ;
SL8_row10(14)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) ;
SL8_row10(15)<=SL8_TS(124) or SL8_TS(125) or SL8_TS(126) or SL8_TS(127) ;
SL8_row10(16)<=SL8_TS(127) or SL8_TS(128) or SL8_TS(129) or SL8_TS(130) ;
SL8_row10(17)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) ;
SL8_row10(18)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) ;
SL8_row10(19)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) ;
SL8_row10(20)<=SL8_TS(136) or SL8_TS(137) or SL8_TS(138) or SL8_TS(139) ;
SL8_row10(21)<=SL8_TS(139) or SL8_TS(140) or SL8_TS(141) or SL8_TS(142) ;
SL8_row10(22)<=SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) ;
SL8_row10(23)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) ;
SL8_row10(24)<=SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) ;
SL8_row10(25)<=SL8_TS(148) or SL8_TS(149) or SL8_TS(150) or SL8_TS(151) ;
SL8_row10(26)<=SL8_TS(151) or SL8_TS(152) or SL8_TS(153) or SL8_TS(154) ;
SL8_row10(27)<=SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) ;
SL8_row10(28)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) ;
SL8_row10(29)<=SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) ;
SL8_row10(30)<=SL8_TS(160) or SL8_TS(161) or SL8_TS(162) or SL8_TS(163) ;
SL8_row10(31)<=SL8_TS(163) or SL8_TS(164) or SL8_TS(165) or SL8_TS(166) ;
SL8_row10(32)<=SL8_TS(165) or SL8_TS(166) or SL8_TS(167) or SL8_TS(168) ;
SL8_row10(33)<=SL8_TS(168) or SL8_TS(169) or SL8_TS(170) ;
SL8_row10(34)<=SL8_TS(170) or SL8_TS(171) or SL8_TS(172) or SL8_TS(173) ;
SL8_row10(35)<=SL8_TS(172) or SL8_TS(173) or SL8_TS(174) or SL8_TS(175) ;
SL8_row10(36)<=SL8_TS(175) or SL8_TS(176) or SL8_TS(177) or SL8_TS(178) ;
SL8_row10(37)<=SL8_TS(177) or SL8_TS(178) or SL8_TS(179) or SL8_TS(180) ;
SL8_row10(38)<=SL8_TS(180) or SL8_TS(181) or SL8_TS(182) ;
SL8_row10(39)<=SL8_TS(182) or SL8_TS(183) or SL8_TS(184) or SL8_TS(185) ;
SL8_row11(0)<=SL8_TS(90) or SL8_TS(91) or SL8_TS(92) ;
SL8_row11(1)<=SL8_TS(92) or SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row11(2)<=SL8_TS(95) or SL8_TS(96) or SL8_TS(97) ;
SL8_row11(3)<=SL8_TS(97) or SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row11(4)<=SL8_TS(99) or SL8_TS(100) or SL8_TS(101) or SL8_TS(102) ;
SL8_row11(5)<=SL8_TS(102) or SL8_TS(103) or SL8_TS(104) ;
SL8_row11(6)<=SL8_TS(104) or SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row11(7)<=SL8_TS(107) or SL8_TS(108) or SL8_TS(109) ;
SL8_row11(8)<=SL8_TS(109) or SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row11(9)<=SL8_TS(111) or SL8_TS(112) or SL8_TS(113) or SL8_TS(114) ;
SL8_row11(10)<=SL8_TS(114) or SL8_TS(115) or SL8_TS(116) ;
SL8_row11(11)<=SL8_TS(116) or SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row11(12)<=SL8_TS(119) or SL8_TS(120) or SL8_TS(121) ;
SL8_row11(13)<=SL8_TS(121) or SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row11(14)<=SL8_TS(123) or SL8_TS(124) or SL8_TS(125) or SL8_TS(126) ;
SL8_row11(15)<=SL8_TS(126) or SL8_TS(127) or SL8_TS(128) ;
SL8_row11(16)<=SL8_TS(128) or SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row11(17)<=SL8_TS(131) or SL8_TS(132) or SL8_TS(133) ;
SL8_row11(18)<=SL8_TS(133) or SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row11(19)<=SL8_TS(135) or SL8_TS(136) or SL8_TS(137) or SL8_TS(138) ;
SL8_row11(20)<=SL8_TS(138) or SL8_TS(139) or SL8_TS(140) ;
SL8_row11(21)<=SL8_TS(140) or SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row11(22)<=SL8_TS(143) or SL8_TS(144) or SL8_TS(145) ;
SL8_row11(23)<=SL8_TS(145) or SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row11(24)<=SL8_TS(147) or SL8_TS(148) or SL8_TS(149) or SL8_TS(150) ;
SL8_row11(25)<=SL8_TS(150) or SL8_TS(151) or SL8_TS(152) ;
SL8_row11(26)<=SL8_TS(152) or SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row11(27)<=SL8_TS(155) or SL8_TS(156) or SL8_TS(157) ;
SL8_row11(28)<=SL8_TS(157) or SL8_TS(158) or SL8_TS(159) or SL8_TS(160) ;
SL8_row11(29)<=SL8_TS(159) or SL8_TS(160) or SL8_TS(161) or SL8_TS(162) ;
SL8_row11(30)<=SL8_TS(162) or SL8_TS(163) or SL8_TS(164) ;
SL8_row11(31)<=SL8_TS(164) or SL8_TS(165) or SL8_TS(166) or SL8_TS(167) ;
SL8_row11(32)<=SL8_TS(167) or SL8_TS(168) or SL8_TS(169) ;
SL8_row11(33)<=SL8_TS(169) or SL8_TS(170) or SL8_TS(171) or SL8_TS(172) ;
SL8_row11(34)<=SL8_TS(171) or SL8_TS(172) or SL8_TS(173) or SL8_TS(174) ;
SL8_row11(35)<=SL8_TS(174) or SL8_TS(175) or SL8_TS(176) ;
SL8_row11(36)<=SL8_TS(176) or SL8_TS(177) or SL8_TS(178) or SL8_TS(179) ;
SL8_row11(37)<=SL8_TS(179) or SL8_TS(180) or SL8_TS(181) ;
SL8_row11(38)<=SL8_TS(181) or SL8_TS(182) or SL8_TS(183) or SL8_TS(184) ;
SL8_row11(39)<=SL8_TS(183) or SL8_TS(184) or SL8_TS(185) or SL8_TS(186) ;
SL8_row12(0)<=SL8_TS(91) or SL8_TS(92) or SL8_TS(93) ;
SL8_row12(1)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) or SL8_TS(96) ;
SL8_row12(2)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) ;
SL8_row12(3)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) or SL8_TS(101) ;
SL8_row12(4)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) ;
SL8_row12(5)<=SL8_TS(103) or SL8_TS(104) or SL8_TS(105) ;
SL8_row12(6)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) or SL8_TS(108) ;
SL8_row12(7)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) ;
SL8_row12(8)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) or SL8_TS(113) ;
SL8_row12(9)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) ;
SL8_row12(10)<=SL8_TS(115) or SL8_TS(116) or SL8_TS(117) ;
SL8_row12(11)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) or SL8_TS(120) ;
SL8_row12(12)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) ;
SL8_row12(13)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) or SL8_TS(125) ;
SL8_row12(14)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) ;
SL8_row12(15)<=SL8_TS(127) or SL8_TS(128) or SL8_TS(129) ;
SL8_row12(16)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) or SL8_TS(132) ;
SL8_row12(17)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) ;
SL8_row12(18)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) or SL8_TS(137) ;
SL8_row12(19)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) ;
SL8_row12(20)<=SL8_TS(139) or SL8_TS(140) or SL8_TS(141) ;
SL8_row12(21)<=SL8_TS(141) or SL8_TS(142) or SL8_TS(143) or SL8_TS(144) ;
SL8_row12(22)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) ;
SL8_row12(23)<=SL8_TS(146) or SL8_TS(147) or SL8_TS(148) or SL8_TS(149) ;
SL8_row12(24)<=SL8_TS(149) or SL8_TS(150) or SL8_TS(151) ;
SL8_row12(25)<=SL8_TS(151) or SL8_TS(152) or SL8_TS(153) ;
SL8_row12(26)<=SL8_TS(153) or SL8_TS(154) or SL8_TS(155) or SL8_TS(156) ;
SL8_row12(27)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) ;
SL8_row12(28)<=SL8_TS(158) or SL8_TS(159) or SL8_TS(160) or SL8_TS(161) ;
SL8_row12(29)<=SL8_TS(161) or SL8_TS(162) or SL8_TS(163) ;
SL8_row12(30)<=SL8_TS(163) or SL8_TS(164) or SL8_TS(165) ;
SL8_row12(31)<=SL8_TS(165) or SL8_TS(166) or SL8_TS(167) or SL8_TS(168) ;
SL8_row12(32)<=SL8_TS(168) or SL8_TS(169) or SL8_TS(170) ;
SL8_row12(33)<=SL8_TS(170) or SL8_TS(171) or SL8_TS(172) or SL8_TS(173) ;
SL8_row12(34)<=SL8_TS(173) or SL8_TS(174) or SL8_TS(175) ;
SL8_row12(35)<=SL8_TS(175) or SL8_TS(176) or SL8_TS(177) ;
SL8_row12(36)<=SL8_TS(177) or SL8_TS(178) or SL8_TS(179) or SL8_TS(180) ;
SL8_row12(37)<=SL8_TS(180) or SL8_TS(181) or SL8_TS(182) ;
SL8_row12(38)<=SL8_TS(182) or SL8_TS(183) or SL8_TS(184) or SL8_TS(185) ;
SL8_row12(39)<=SL8_TS(185) or SL8_TS(186) or SL8_TS(187) ;
SL8_row13(0)<=SL8_TS(92) or SL8_TS(93) or SL8_TS(94) ;
SL8_row13(1)<=SL8_TS(94) or SL8_TS(95) or SL8_TS(96) or SL8_TS(97) ;
SL8_row13(2)<=SL8_TS(97) or SL8_TS(98) or SL8_TS(99) ;
SL8_row13(3)<=SL8_TS(99) or SL8_TS(100) or SL8_TS(101) ;
SL8_row13(4)<=SL8_TS(102) or SL8_TS(103) or SL8_TS(104) ;
SL8_row13(5)<=SL8_TS(104) or SL8_TS(105) or SL8_TS(106) ;
SL8_row13(6)<=SL8_TS(106) or SL8_TS(107) or SL8_TS(108) or SL8_TS(109) ;
SL8_row13(7)<=SL8_TS(109) or SL8_TS(110) or SL8_TS(111) ;
SL8_row13(8)<=SL8_TS(111) or SL8_TS(112) or SL8_TS(113) ;
SL8_row13(9)<=SL8_TS(114) or SL8_TS(115) or SL8_TS(116) ;
SL8_row13(10)<=SL8_TS(116) or SL8_TS(117) or SL8_TS(118) ;
SL8_row13(11)<=SL8_TS(118) or SL8_TS(119) or SL8_TS(120) or SL8_TS(121) ;
SL8_row13(12)<=SL8_TS(121) or SL8_TS(122) or SL8_TS(123) ;
SL8_row13(13)<=SL8_TS(123) or SL8_TS(124) or SL8_TS(125) ;
SL8_row13(14)<=SL8_TS(126) or SL8_TS(127) or SL8_TS(128) ;
SL8_row13(15)<=SL8_TS(128) or SL8_TS(129) or SL8_TS(130) ;
SL8_row13(16)<=SL8_TS(130) or SL8_TS(131) or SL8_TS(132) or SL8_TS(133) ;
SL8_row13(17)<=SL8_TS(133) or SL8_TS(134) or SL8_TS(135) ;
SL8_row13(18)<=SL8_TS(135) or SL8_TS(136) or SL8_TS(137) ;
SL8_row13(19)<=SL8_TS(138) or SL8_TS(139) or SL8_TS(140) ;
SL8_row13(20)<=SL8_TS(140) or SL8_TS(141) or SL8_TS(142) ;
SL8_row13(21)<=SL8_TS(142) or SL8_TS(143) or SL8_TS(144) or SL8_TS(145) ;
SL8_row13(22)<=SL8_TS(145) or SL8_TS(146) or SL8_TS(147) ;
SL8_row13(23)<=SL8_TS(147) or SL8_TS(148) or SL8_TS(149) ;
SL8_row13(24)<=SL8_TS(150) or SL8_TS(151) or SL8_TS(152) ;
SL8_row13(25)<=SL8_TS(152) or SL8_TS(153) or SL8_TS(154) ;
SL8_row13(26)<=SL8_TS(154) or SL8_TS(155) or SL8_TS(156) or SL8_TS(157) ;
SL8_row13(27)<=SL8_TS(157) or SL8_TS(158) or SL8_TS(159) ;
SL8_row13(28)<=SL8_TS(159) or SL8_TS(160) or SL8_TS(161) ;
SL8_row13(29)<=SL8_TS(162) or SL8_TS(163) or SL8_TS(164) ;
SL8_row13(30)<=SL8_TS(164) or SL8_TS(165) or SL8_TS(166) ;
SL8_row13(31)<=SL8_TS(166) or SL8_TS(167) or SL8_TS(168) or SL8_TS(169) ;
SL8_row13(32)<=SL8_TS(169) or SL8_TS(170) or SL8_TS(171) ;
SL8_row13(33)<=SL8_TS(171) or SL8_TS(172) or SL8_TS(173) ;
SL8_row13(34)<=SL8_TS(174) or SL8_TS(175) or SL8_TS(176) ;
SL8_row13(35)<=SL8_TS(176) or SL8_TS(177) or SL8_TS(178) ;
SL8_row13(36)<=SL8_TS(178) or SL8_TS(179) or SL8_TS(180) or SL8_TS(181) ;
SL8_row13(37)<=SL8_TS(181) or SL8_TS(182) or SL8_TS(183) ;
SL8_row13(38)<=SL8_TS(183) or SL8_TS(184) or SL8_TS(185) ;
SL8_row13(39)<=SL8_TS(186) or SL8_TS(187) or SL8_TS(188) ;
SL8_row14(0)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row14(1)<=SL8_TS(95) or SL8_TS(96) or SL8_TS(97) ;
SL8_row14(2)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row14(3)<=SL8_TS(100) or SL8_TS(101) or SL8_TS(102) ;
SL8_row14(4)<=SL8_TS(102) or SL8_TS(103) or SL8_TS(104) ;
SL8_row14(5)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row14(6)<=SL8_TS(107) or SL8_TS(108) or SL8_TS(109) ;
SL8_row14(7)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row14(8)<=SL8_TS(112) or SL8_TS(113) or SL8_TS(114) ;
SL8_row14(9)<=SL8_TS(114) or SL8_TS(115) or SL8_TS(116) ;
SL8_row14(10)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row14(11)<=SL8_TS(119) or SL8_TS(120) or SL8_TS(121) ;
SL8_row14(12)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row14(13)<=SL8_TS(124) or SL8_TS(125) or SL8_TS(126) ;
SL8_row14(14)<=SL8_TS(126) or SL8_TS(127) or SL8_TS(128) ;
SL8_row14(15)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row14(16)<=SL8_TS(131) or SL8_TS(132) or SL8_TS(133) ;
SL8_row14(17)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row14(18)<=SL8_TS(136) or SL8_TS(137) or SL8_TS(138) ;
SL8_row14(19)<=SL8_TS(138) or SL8_TS(139) or SL8_TS(140) ;
SL8_row14(20)<=SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row14(21)<=SL8_TS(143) or SL8_TS(144) or SL8_TS(145) ;
SL8_row14(22)<=SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row14(23)<=SL8_TS(148) or SL8_TS(149) or SL8_TS(150) ;
SL8_row14(24)<=SL8_TS(150) or SL8_TS(151) or SL8_TS(152) ;
SL8_row14(25)<=SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row14(26)<=SL8_TS(155) or SL8_TS(156) or SL8_TS(157) ;
SL8_row14(27)<=SL8_TS(158) or SL8_TS(159) or SL8_TS(160) ;
SL8_row14(28)<=SL8_TS(160) or SL8_TS(161) or SL8_TS(162) ;
SL8_row14(29)<=SL8_TS(162) or SL8_TS(163) or SL8_TS(164) ;
SL8_row14(30)<=SL8_TS(165) or SL8_TS(166) or SL8_TS(167) ;
SL8_row14(31)<=SL8_TS(167) or SL8_TS(168) or SL8_TS(169) ;
SL8_row14(32)<=SL8_TS(170) or SL8_TS(171) or SL8_TS(172) ;
SL8_row14(33)<=SL8_TS(172) or SL8_TS(173) or SL8_TS(174) ;
SL8_row14(34)<=SL8_TS(174) or SL8_TS(175) or SL8_TS(176) ;
SL8_row14(35)<=SL8_TS(177) or SL8_TS(178) or SL8_TS(179) ;
SL8_row14(36)<=SL8_TS(179) or SL8_TS(180) or SL8_TS(181) ;
SL8_row14(37)<=SL8_TS(182) or SL8_TS(183) or SL8_TS(184) ;
SL8_row14(38)<=SL8_TS(184) or SL8_TS(185) or SL8_TS(186) ;
SL8_row14(39)<=SL8_TS(186) or SL8_TS(187) or SL8_TS(188) ;
SL8_row15(0)<=SL8_TS(93) or SL8_TS(94) or SL8_TS(95) ;
SL8_row15(1)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) ;
SL8_row15(2)<=SL8_TS(98) or SL8_TS(99) or SL8_TS(100) ;
SL8_row15(3)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) ;
SL8_row15(4)<=SL8_TS(103) or SL8_TS(104) or SL8_TS(105) ;
SL8_row15(5)<=SL8_TS(105) or SL8_TS(106) or SL8_TS(107) ;
SL8_row15(6)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) ;
SL8_row15(7)<=SL8_TS(110) or SL8_TS(111) or SL8_TS(112) ;
SL8_row15(8)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) ;
SL8_row15(9)<=SL8_TS(115) or SL8_TS(116) or SL8_TS(117) ;
SL8_row15(10)<=SL8_TS(117) or SL8_TS(118) or SL8_TS(119) ;
SL8_row15(11)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) ;
SL8_row15(12)<=SL8_TS(122) or SL8_TS(123) or SL8_TS(124) ;
SL8_row15(13)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) ;
SL8_row15(14)<=SL8_TS(127) or SL8_TS(128) or SL8_TS(129) ;
SL8_row15(15)<=SL8_TS(129) or SL8_TS(130) or SL8_TS(131) ;
SL8_row15(16)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) ;
SL8_row15(17)<=SL8_TS(134) or SL8_TS(135) or SL8_TS(136) ;
SL8_row15(18)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) ;
SL8_row15(19)<=SL8_TS(139) or SL8_TS(140) or SL8_TS(141) ;
SL8_row15(20)<=SL8_TS(141) or SL8_TS(142) or SL8_TS(143) ;
SL8_row15(21)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) ;
SL8_row15(22)<=SL8_TS(146) or SL8_TS(147) or SL8_TS(148) ;
SL8_row15(23)<=SL8_TS(149) or SL8_TS(150) or SL8_TS(151) ;
SL8_row15(24)<=SL8_TS(151) or SL8_TS(152) or SL8_TS(153) ;
SL8_row15(25)<=SL8_TS(153) or SL8_TS(154) or SL8_TS(155) ;
SL8_row15(26)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) ;
SL8_row15(27)<=SL8_TS(158) or SL8_TS(159) or SL8_TS(160) ;
SL8_row15(28)<=SL8_TS(161) or SL8_TS(162) or SL8_TS(163) ;
SL8_row15(29)<=SL8_TS(163) or SL8_TS(164) or SL8_TS(165) ;
SL8_row15(30)<=SL8_TS(165) or SL8_TS(166) or SL8_TS(167) ;
SL8_row15(31)<=SL8_TS(168) or SL8_TS(169) or SL8_TS(170) ;
SL8_row15(32)<=SL8_TS(170) or SL8_TS(171) or SL8_TS(172) ;
SL8_row15(33)<=SL8_TS(173) or SL8_TS(174) or SL8_TS(175) ;
SL8_row15(34)<=SL8_TS(175) or SL8_TS(176) or SL8_TS(177) ;
SL8_row15(35)<=SL8_TS(177) or SL8_TS(178) or SL8_TS(179) ;
SL8_row15(36)<=SL8_TS(180) or SL8_TS(181) or SL8_TS(182) ;
SL8_row15(37)<=SL8_TS(182) or SL8_TS(183) or SL8_TS(184) ;
SL8_row15(38)<=SL8_TS(185) or SL8_TS(186) or SL8_TS(187) ;
SL8_row15(39)<=SL8_TS(187) or SL8_TS(188) or SL8_TS(189) ;
SL8_row16(0)<=SL8_TS(94) or SL8_TS(95) or SL8_TS(96) ;
SL8_row16(1)<=SL8_TS(96) or SL8_TS(97) or SL8_TS(98) ;
SL8_row16(2)<=SL8_TS(99) or SL8_TS(100) or SL8_TS(101) ;
SL8_row16(3)<=SL8_TS(101) or SL8_TS(102) or SL8_TS(103) ;
SL8_row16(4)<=SL8_TS(104) or SL8_TS(105) ;
SL8_row16(5)<=SL8_TS(106) or SL8_TS(107) or SL8_TS(108) ;
SL8_row16(6)<=SL8_TS(108) or SL8_TS(109) or SL8_TS(110) ;
SL8_row16(7)<=SL8_TS(111) or SL8_TS(112) or SL8_TS(113) ;
SL8_row16(8)<=SL8_TS(113) or SL8_TS(114) or SL8_TS(115) ;
SL8_row16(9)<=SL8_TS(116) or SL8_TS(117) ;
SL8_row16(10)<=SL8_TS(118) or SL8_TS(119) or SL8_TS(120) ;
SL8_row16(11)<=SL8_TS(120) or SL8_TS(121) or SL8_TS(122) ;
SL8_row16(12)<=SL8_TS(123) or SL8_TS(124) or SL8_TS(125) ;
SL8_row16(13)<=SL8_TS(125) or SL8_TS(126) or SL8_TS(127) ;
SL8_row16(14)<=SL8_TS(128) or SL8_TS(129) ;
SL8_row16(15)<=SL8_TS(130) or SL8_TS(131) or SL8_TS(132) ;
SL8_row16(16)<=SL8_TS(132) or SL8_TS(133) or SL8_TS(134) ;
SL8_row16(17)<=SL8_TS(135) or SL8_TS(136) or SL8_TS(137) ;
SL8_row16(18)<=SL8_TS(137) or SL8_TS(138) or SL8_TS(139) ;
SL8_row16(19)<=SL8_TS(140) or SL8_TS(141) ;
SL8_row16(20)<=SL8_TS(142) or SL8_TS(143) or SL8_TS(144) ;
SL8_row16(21)<=SL8_TS(144) or SL8_TS(145) or SL8_TS(146) ;
SL8_row16(22)<=SL8_TS(147) or SL8_TS(148) or SL8_TS(149) ;
SL8_row16(23)<=SL8_TS(149) or SL8_TS(150) or SL8_TS(151) ;
SL8_row16(24)<=SL8_TS(152) or SL8_TS(153) ;
SL8_row16(25)<=SL8_TS(154) or SL8_TS(155) or SL8_TS(156) ;
SL8_row16(26)<=SL8_TS(156) or SL8_TS(157) or SL8_TS(158) ;
SL8_row16(27)<=SL8_TS(159) or SL8_TS(160) or SL8_TS(161) ;
SL8_row16(28)<=SL8_TS(161) or SL8_TS(162) or SL8_TS(163) ;
SL8_row16(29)<=SL8_TS(164) or SL8_TS(165) ;
SL8_row16(30)<=SL8_TS(166) or SL8_TS(167) or SL8_TS(168) ;
SL8_row16(31)<=SL8_TS(168) or SL8_TS(169) or SL8_TS(170) ;
SL8_row16(32)<=SL8_TS(171) or SL8_TS(172) or SL8_TS(173) ;
SL8_row16(33)<=SL8_TS(173) or SL8_TS(174) or SL8_TS(175) ;
SL8_row16(34)<=SL8_TS(176) or SL8_TS(177) ;
SL8_row16(35)<=SL8_TS(178) or SL8_TS(179) or SL8_TS(180) ;
SL8_row16(36)<=SL8_TS(180) or SL8_TS(181) or SL8_TS(182) ;
SL8_row16(37)<=SL8_TS(183) or SL8_TS(184) or SL8_TS(185) ;
SL8_row16(38)<=SL8_TS(185) or SL8_TS(186) or SL8_TS(187) ;
SL8_row16(39)<=SL8_TS(188) or SL8_TS(189) ;
 
end Behavioral;
